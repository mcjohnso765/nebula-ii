* NGSPICE file created from team_02_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_02_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_185_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_176_Left_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] net896 net943 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11834__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ net73 team_02_WB.START_ADDR_VAL_REG\[10\] net956 vssd1 vssd1 vccd1 vccd1
+ _02638_ sky130_fd_sc_hd__mux2_1
XANTENNA__11618__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _04214_ _04215_ net651 net792 net1518 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08484_ _03321_ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12665__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_185_Left_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13350__A team_02_WB.instance_to_wrap.ramload\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] net709 _04616_ _04618_
+ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10038__X _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09036_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\] net924 net920 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout796_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold340 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10357__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_X net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 team_02_WB.instance_to_wrap.top.a1.row1\[56\] vssd1 vssd1 vccd1 vccd1 net1724
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09762__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _04514_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08970__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 _04508_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_4
X_09938_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\] net816 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\]
+ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a221o_1
Xfanout842 _04400_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_8
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_2
Xfanout864 _04543_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_8
Xfanout875 _04539_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09514__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 net889 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_8
X_09869_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\] net737 net677 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\]
+ _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a221o_1
Xfanout897 _04531_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1040 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11744__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net345 net2083 net487 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__mux2_1
Xhold1073 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _07387_ _07399_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__nand2_1
Xhold1084 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ net339 net1856 net588 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10587__C _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14550_ net1106 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
X_11762_ net335 net1792 net599 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13501_ net2586 _04268_ _04346_ team_02_WB.instance_to_wrap.top.ru.next_read_i vssd1
+ vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__o31a_1
X_10713_ team_02_WB.instance_to_wrap.top.pc\[22\] _06177_ _06229_ vssd1 vssd1 vccd1
+ vccd1 _06230_ sky130_fd_sc_hd__a21o_1
X_14481_ net1233 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XANTENNA__12575__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10884__A _06080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ _07138_ _07174_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__a21o_1
XANTENNA__11332__X _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16725__1280 vssd1 vssd1 vccd1 vccd1 _16725__1280/HI net1280 sky130_fd_sc_hd__conb_1
X_16220_ clknet_leaf_20_wb_clk_i _02360_ _01028_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input92_A wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] _03023_ _03039_ vssd1
+ vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__o21ai_2
X_10644_ _04338_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16151_ clknet_leaf_120_wb_clk_i _02291_ _00959_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10575_ net528 net406 _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ net1590 net1018 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[25\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_106_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold796_X net2158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15102_ net1081 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XANTENNA__10060__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ net250 net2012 net566 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__mux2_1
X_16082_ clknet_leaf_76_wb_clk_i _02222_ _00890_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13294_ net1631 net985 net964 _02996_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15033_ net1228 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
XANTENNA__11919__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ net245 net2436 net573 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__mux2_1
XANTENNA__10348__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14091__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ net349 net1912 net462 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08961__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15935_ clknet_leaf_60_wb_clk_i _02075_ _00743_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11058_ _06431_ _06433_ net393 vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__mux2_1
XANTENNA__09505__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11312__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] net780 net719 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_199_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15866_ clknet_leaf_19_wb_clk_i _02006_ _00674_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08529__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14817_ net1256 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15797_ clknet_leaf_31_wb_clk_i _01937_ _00605_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14748_ net1194 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12485__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14679_ net1219 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07579__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16418_ clknet_leaf_80_wb_clk_i _02553_ _01226_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16349_ clknet_leaf_12_wb_clk_i _02489_ _01157_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09647__X _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11829__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07984_ _03601_ _03662_ _03675_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__mux2_1
X_09723_ _05233_ _05235_ _05237_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13345__A team_02_WB.instance_to_wrap.ramload\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09654_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\] net788 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a22o_1
XANTENNA__08439__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08605_ net91 net1536 net956 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\] net745 _05097_ _05098_
+ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_fanout544_A _04498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08536_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\] _04177_ vssd1 vssd1 vccd1
+ vccd1 _04221_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_193_Left_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net1578 net1006 net981 _04167_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12395__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_A _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08398_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_4
Xwire517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
XFILLER_0_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_4
XFILLER_0_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1241_X net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10360_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__inv_2
XANTENNA__09983__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11739__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09019_ _04297_ net944 _04509_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10291_ _05788_ net619 net968 vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__mux2_1
X_12030_ net319 net2048 net474 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold170 team_02_WB.START_ADDR_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold192 _02614_ vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout650 _04331_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
Xfanout672 _04469_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
X_13981_ net1204 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
Xfanout683 _04402_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_6
Xfanout694 _04394_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_4
XANTENNA__13295__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ clknet_leaf_25_wb_clk_i _01860_ _00528_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12932_ team_02_WB.instance_to_wrap.top.pc\[26\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _07452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ clknet_leaf_9_wb_clk_i _01791_ _00459_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12863_ _07381_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13047__A2 _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14602_ net1189 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
X_11814_ net269 net2626 net589 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
X_15582_ clknet_leaf_3_wb_clk_i _01722_ _00390_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12794_ net378 _06534_ _07076_ _07127_ _06037_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_194_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09120__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ net1114 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
X_11745_ net265 net2180 net598 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10281__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14464_ net1105 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
X_11676_ _05187_ _05206_ _05979_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16203_ clknet_leaf_16_wb_clk_i _02343_ _01011_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13415_ _03018_ _03024_ _03025_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_64_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10627_ team_02_WB.instance_to_wrap.top.pc\[27\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _06144_ sky130_fd_sc_hd__nor2_1
X_14395_ net1076 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10033__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16134_ clknet_leaf_9_wb_clk_i _02274_ _00942_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13346_ team_02_WB.instance_to_wrap.ramload\[8\] net1015 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[8\] sky130_fd_sc_hd__and2_1
X_10558_ _04755_ net387 vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10553__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16065_ clknet_leaf_100_wb_clk_i _02205_ _00873_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13277_ team_02_WB.instance_to_wrap.top.pc\[21\] net1053 _06679_ net935 vssd1 vssd1
+ vccd1 vccd1 _02988_ sky130_fd_sc_hd__a22o_1
X_10489_ _05919_ _06005_ _05920_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_121_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09187__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15016_ net1146 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XANTENNA__09726__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net1715 net296 net614 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ net295 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\] net464 vssd1
+ vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
XANTENNA__10789__A _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16412__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15918_ clknet_leaf_45_wb_clk_i _02058_ _00726_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire512_A _05488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15849_ clknet_leaf_115_wb_clk_i _01989_ _00657_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09370_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] net896 net943 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ _04028_ _04032_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08706__B _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ _03957_ _03960_ _03945_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10272__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _03882_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_41_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09818__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09965__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput220 net220 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03687_ _03688_ vssd1 vssd1
+ vccd1 vccd1 _03690_ sky130_fd_sc_hd__or3_1
XANTENNA__13277__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\] net698 _05219_ _05220_
+ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a2111o_1
X_07898_ _03591_ _03620_ net316 vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__o21a_1
XANTENNA__09350__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09637_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\] net864 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout926_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\] net722 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\]
+ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08519_ team_02_WB.instance_to_wrap.top.a1.data\[4\] net958 vssd1 vssd1 vccd1 vccd1
+ _04208_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ _05009_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_176_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11530_ _06037_ net384 _06296_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__a31oi_2
XANTENNA__10263__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ _05512_ _05514_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__nand2_2
XFILLER_0_162_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ net1019 _02953_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__or2_1
XANTENNA__10015__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ _05465_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__or2_1
X_14180_ net1136 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XANTENNA__09956__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11392_ net604 _06884_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__and3_2
XFILLER_0_104_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10566__A3 _06080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ _06887_ net232 _02898_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__o22a_1
X_10343_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\] net721 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a22o_1
XANTENNA__09708__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\] net828 net816 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\]
+ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a221o_1
XANTENNA_input55_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _07455_ _07456_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_72_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15238__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net253 net2253 net477 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_6
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout491 _07196_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
X_16752_ net1296 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XANTENNA__11279__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11279__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13964_ net1244 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XANTENNA_input10_X net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ clknet_leaf_120_wb_clk_i _01843_ _00511_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12915_ _07359_ _07434_ _07358_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__a21oi_1
X_16683_ clknet_leaf_65_wb_clk_i _02800_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11304__A1_N net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13895_ net1244 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XANTENNA__11932__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15634_ clknet_leaf_54_wb_clk_i _01774_ _00442_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ _05061_ _06186_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15565_ clknet_leaf_48_wb_clk_i _01705_ _00373_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12777_ _06548_ _06674_ _07266_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_83_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14516_ net1238 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
X_11728_ net336 net2620 net603 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XANTENNA__10254__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15496_ clknet_leaf_11_wb_clk_i _01636_ _00304_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14447_ net1197 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _05832_ _05910_ _06429_ _07142_ _07144_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_211_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11520__X _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11203__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14378_ net1117 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold906 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ clknet_leaf_31_wb_clk_i _02257_ _00925_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16532__Q team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold917 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap636 _04564_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_2
X_13329_ team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] team_02_WB.instance_to_wrap.top.a1.nextHex\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[0\] sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_114_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold928 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 team_02_WB.instance_to_wrap.top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 net2301
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16048_ clknet_leaf_23_wb_clk_i _02188_ _00856_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08870_ net1057 net1032 team_02_WB.instance_to_wrap.wb.prev_BUSY_O vssd1 vssd1 vccd1
+ vccd1 _04432_ sky130_fd_sc_hd__or3b_4
XFILLER_0_208_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_209_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07821_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] _03541_ _03542_ vssd1 vssd1
+ vccd1 vccd1 _03544_ sky130_fd_sc_hd__or3_1
XFILLER_0_208_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12003__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _03461_ _03462_ _03453_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a21o_1
XANTENNA__09332__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07683_ _03375_ _03404_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11842__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09422_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\] net892 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07621__A team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09353_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] net780 _04868_ _04869_
+ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a211o_1
XANTENNA__08438__A2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13431__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08304_ net2301 net1007 net980 _04018_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10245__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09284_ _04794_ _04796_ _04798_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nor4_2
XFILLER_0_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ _03950_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12673__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1151_A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09938__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ _03839_ _03859_ _03838_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11289__S net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08097_ net1662 net1007 net980 _03817_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload90 clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_8
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09571__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ net1058 _04499_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__or4bb_4
XANTENNA__13236__C _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_117_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ _06078_ _06100_ net407 vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_206_Right_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12700_ net359 net1784 net433 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__mux2_1
X_13680_ _03206_ _03210_ net1141 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a21oi_1
X_10892_ net380 _06404_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ net1681 net330 net552 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10236__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15350_ clknet_leaf_57_wb_clk_i _01490_ _00163_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_183_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ net323 net1702 net443 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ net1181 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
X_11513_ net668 _06995_ _06996_ net836 _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__o221a_1
XANTENNA__12583__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ clknet_leaf_70_wb_clk_i _01425_ _00094_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ net305 net2502 net559 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14232_ net1189 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
X_11444_ _06848_ _06939_ net397 vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__mux2_1
XANTENNA__09929__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14163_ net1078 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
X_11375_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_189_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ net976 _07420_ _02882_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o31ai_1
X_10326_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] net820 net914 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a22o_1
X_14094_ net1082 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15195__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11927__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13045_ _07436_ _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__xor2_1
X_10257_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\] net718 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a22o_1
XANTENNA__10942__A2_N net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1220 net1223 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1231 net1236 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_4
X_10188_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\] net815 net913 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\]
+ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a221o_1
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__buf_4
Xfanout1253 net1255 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_4
Xfanout1264 net1265 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_4_14__f_wb_clk_i_X clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14996_ net1133 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XANTENNA__09314__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16735_ net1281 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_0_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13947_ net1243 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14539__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16666_ clknet_leaf_70_wb_clk_i _02785_ _01408_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13878_ net1253 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15617_ clknet_leaf_101_wb_clk_i _01757_ _00425_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ team_02_WB.instance_to_wrap.top.i_ready team_02_WB.instance_to_wrap.top.testpc.en_latched
+ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__nand2b_2
X_16597_ clknet_leaf_89_wb_clk_i _02716_ _01390_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10227__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15548_ clknet_leaf_20_wb_clk_i _01688_ _00356_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12493__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15479_ clknet_leaf_120_wb_clk_i _01619_ _00287_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_08020_ _03733_ _03737_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold703 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold769 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\] net726 _05470_ _05482_
+ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11837__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ net1436 _04443_ net930 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08853_ net141 net1039 net1037 net1496 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07804_ _03481_ _03513_ _03526_ _03485_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a22o_1
X_08784_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] net777 net749 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a22o_1
XANTENNA__13637__C1 _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09305__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13101__B2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ _03420_ _03427_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__and2_1
XANTENNA__12668__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout457_A _07221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08718__Y _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1199_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13353__A team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07666_ _03356_ _03360_ _03357_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_140_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09405_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\] net782 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__a22o_1
X_07597_ net1749 net1008 net980 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09336_ _04846_ _04848_ _04850_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or4_1
XANTENNA__10218__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\] net775 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _03918_ _03927_ _03917_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__and3b_1
XANTENNA__13168__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09198_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] net895 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08149_ _03863_ _03866_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09792__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ net423 _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11747__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\] net824 net821 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a22o_1
X_11091_ _05972_ _06023_ _06597_ _05975_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o22a_1
XANTENNA__09284__Y _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__nand2_2
XANTENNA__12789__D _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 team_02_WB.instance_to_wrap.ramstore\[12\] vssd1 vssd1 vccd1 vccd1 net1392
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 _02620_ vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold52 team_02_WB.START_ADDR_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1129 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold63 _02602_ vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_02_WB.instance_to_wrap.top.a1.data\[3\] vssd1 vssd1 vccd1 vccd1 net1436
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 _02600_ vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] _03284_
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\] vssd1 vssd1 vccd1
+ vccd1 _03287_ sky130_fd_sc_hd__a21o_1
Xhold96 _02598_ vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ net1203 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12578__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10887__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net298 net2228 net479 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
X_16520_ clknet_leaf_5_wb_clk_i _02654_ _01327_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13732_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] _03240_ vssd1 vssd1 vccd1
+ vccd1 _03242_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10944_ net837 _06426_ _06454_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16451_ clknet_leaf_64_wb_clk_i _02586_ _01259_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13663_ net1367 _04086_ net850 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
X_10875_ net370 _06099_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ clknet_leaf_36_wb_clk_i _01542_ _00210_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12614_ net1990 net263 net553 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__mux2_1
XANTENNA__10209__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16382_ clknet_leaf_88_wb_clk_i _02517_ _01190_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ _03141_ _03144_ _03146_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__or4_1
XFILLER_0_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_85_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15333_ clknet_leaf_43_wb_clk_i _01476_ _00146_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12545_ net250 net2219 net445 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10090__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15264_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[23\]
+ _00077_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_12476_ net247 net2331 net558 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14215_ net1173 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
X_11427_ _06922_ _06923_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__or2_1
XANTENNA_5 _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ net1263 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09783__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14146_ net1129 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ net954 _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__nand2_1
X_10309_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\] net709 _05822_ _05823_
+ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a2111o_1
X_14077_ net1204 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_169_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ net1674 net293 net638 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09535__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ _07545_ _07546_ net230 vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_206_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1050 team_02_WB.instance_to_wrap.top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1
+ net1050 sky130_fd_sc_hd__buf_1
Xfanout1061 team_02_WB.instance_to_wrap.top.a1.instruction\[12\] vssd1 vssd1 vccd1
+ vccd1 net1061 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_177_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1072 net1074 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_4
Xfanout1083 net1085 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_4
XFILLER_0_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1094 net1101 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12488__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1156 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XANTENNA__11245__X _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13173__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16718_ net1350 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_202_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16649_ clknet_leaf_92_wb_clk_i _02768_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09066__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\] net914 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09369__Y _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12076__X _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11421__A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ _04566_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nor2_2
X_08003_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03723_ _03724_ _03722_ vssd1
+ vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__o211a_1
Xhold500 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold533 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold544 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08730__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] net722 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold599 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1114_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ net1522 _04434_ net930 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__a22o_1
Xhold1200 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ net159 net1043 net1035 net1443 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
Xhold1222 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1255 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\] net785 net733 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\]
+ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a221o_1
XANTENNA__12398__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13625__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15520__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07718_ _03402_ _03429_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08698_ net1001 net848 vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__nand2_1
XANTENNA__08501__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ _03370_ _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nor2_1
XANTENNA__14907__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10660_ _06128_ _06176_ _04490_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09057__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15670__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09319_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] net780 net764 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\]
+ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ net380 _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10072__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ net317 net2614 net564 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ net297 net1885 net574 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__mux2_1
X_14000_ net1234 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11212_ net413 _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__nand2_1
XANTENNA__09765__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08640__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ net293 net1781 net577 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__mux2_1
X_11143_ _06229_ _06650_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__nor2_1
XANTENNA__13258__A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13313__B2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15951_ clknet_leaf_41_wb_clk_i _02091_ _00759_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11074_ _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\] net811 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\]
+ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__a221o_1
X_14902_ net1120 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
X_15882_ clknet_leaf_37_wb_clk_i _02022_ _00690_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08639__X _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14833_ net1223 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14764_ net1217 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_201_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12101__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ net242 net2581 net479 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09296__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13715_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] _03231_ net1139 vssd1
+ vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a21oi_1
X_16503_ clknet_leaf_27_wb_clk_i _02637_ _01310_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ _06439_ _06440_ net393 vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14695_ net1180 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
X_16434_ clknet_leaf_44_wb_clk_i net1471 _01242_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dfrtp_1
X_13646_ _03109_ _03113_ net1144 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21o_1
X_10858_ _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand2_2
XANTENNA__09048__A2 _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16365_ clknet_leaf_49_wb_clk_i _02505_ _01173_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13577_ _03106_ net963 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__nand2b_1
X_10789_ _05356_ net404 vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15316_ clknet_leaf_62_wb_clk_i _01459_ _00129_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12528_ net319 net2235 net446 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
X_16296_ clknet_leaf_24_wb_clk_i _02436_ _01104_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10128__Y _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15247_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[6\]
+ _00060_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12459_ net296 net2524 net453 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09756__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15178_ net1142 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09220__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14129_ net1232 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XANTENNA__10291__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 _06840_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09508__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__B2 _03001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09670_ net520 vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ net74 net1495 net955 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12011__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ _04211_ _04212_ net651 net792 net1561 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a32o_1
XANTENNA__11618__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09287__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08483_ net1010 _04168_ net1048 _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11850__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09039__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout322_A _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09104_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\] net693 _04619_ _04620_
+ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] net797 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a22o_1
XANTENNA__12681__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1231_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10990__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold352 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_8
Xfanout821 _04514_ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
X_09937_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\] net906 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a22o_1
Xfanout832 _04506_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
Xfanout843 _04400_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _04559_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_6
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 _04543_ vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_181_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout876 _04539_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_8
X_09868_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] net773 net769 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__a22o_1
Xfanout887 net889 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_8
Xhold1030 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 _04526_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_4
Xhold1041 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ net1607 net1038 net990 team_02_WB.instance_to_wrap.ramaddr\[12\] vssd1 vssd1
+ vccd1 vccd1 _02606_ sky130_fd_sc_hd__a22o_1
Xhold1063 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\] net924 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__a22o_1
Xhold1074 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net332 net2246 net591 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
Xhold1096 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09278__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net325 net1718 net597 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11760__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ net1018 team_02_WB.instance_to_wrap.top.ru.next_dready vssd1 vssd1 vccd1
+ vccd1 _00005_ sky130_fd_sc_hd__or2_1
XANTENNA__10293__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ _06178_ _06228_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__and2_1
X_14480_ net1232 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11692_ _04461_ _06109_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__or3b_1
XFILLER_0_138_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13431_ team_02_WB.instance_to_wrap.top.lcd.currentState\[5\] net962 net1066 vssd1
+ vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10643_ net1001 _06156_ _06158_ _06159_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__or4b_1
XANTENNA__13231__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ clknet_leaf_22_wb_clk_i _02290_ _00958_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input85_A wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ net1696 net1018 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[24\]
+ sky130_fd_sc_hd__and2_1
X_10574_ _05061_ net406 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11793__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ net1104 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12313_ net254 net2146 net565 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16081_ clknet_leaf_128_wb_clk_i _02221_ _00889_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12591__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ _06883_ _02959_ team_02_WB.instance_to_wrap.top.pc\[13\] net1054 vssd1 vssd1
+ vccd1 vccd1 _02996_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14372__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ net1168 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XANTENNA__09738__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ net242 net2287 net573 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09202__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ net351 net1750 net462 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ _06632_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13298__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ net408 _06429_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or2_1
X_15934_ clknet_leaf_1_wb_clk_i _02074_ _00742_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10008_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\] net764 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a22o_1
XANTENNA__09910__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ clknet_leaf_121_wb_clk_i _02005_ _00673_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14816_ net1104 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15796_ clknet_leaf_3_wb_clk_i _01936_ _00604_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09269__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14747_ net1084 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
X_11959_ net298 net2402 net586 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__mux2_1
XANTENNA__10284__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14678_ net1096 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13629_ _03023_ _03106_ _03169_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__or4_1
X_16417_ clknet_leaf_85_wb_clk_i _02552_ _01225_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13222__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10036__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09977__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16348_ clknet_leaf_17_wb_clk_i _02488_ _01156_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08832__X _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09441__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ clknet_leaf_120_wb_clk_i _02419_ _01087_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09729__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10339__A1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13101__A1_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16491__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07983_ _03677_ _03704_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__xor2_1
XANTENNA__13289__B1 _06830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] net821 net883 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\]
+ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a221o_1
X_09653_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\] net719 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a22o_1
X_08604_ net92 net1551 net956 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XANTENNA__11146__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] net673 _05099_ _05100_
+ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ team_02_WB.instance_to_wrap.top.a1.data\[0\] net959 vssd1 vssd1 vccd1 vccd1
+ _04220_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12676__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10275__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13361__A net2514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ _04164_ _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09680__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08483__A3 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13213__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout704_A _04389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _04092_ _04099_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_162_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10027__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire518 _05400_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_2
XFILLER_0_107_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09968__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire529 net531 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08742__X _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10924__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09018_ _04504_ _04519_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__nor2_2
X_10290_ net619 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold160 team_02_WB.instance_to_wrap.top.a1.data\[11\] vssd1 vssd1 vccd1 vccd1 net1522
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 team_02_WB.instance_to_wrap.ramload\[14\] vssd1 vssd1 vccd1 vccd1 net1533
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_02_WB.instance_to_wrap.top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1
+ net1544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold193 team_02_WB.START_ADDR_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _04454_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_4
Xfanout651 _04224_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_2
XANTENNA__11755__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 _06112_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_148_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13980_ net1201 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
Xfanout673 net676 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_4
Xfanout684 _04402_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout695 _04394_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_8
X_12931_ team_02_WB.instance_to_wrap.top.pc\[27\] _06147_ vssd1 vssd1 vccd1 vccd1
+ _07451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ clknet_leaf_118_wb_clk_i _01790_ _00458_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12862_ net515 _05444_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14601_ net1228 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11813_ net261 net2105 net589 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
X_15581_ clknet_leaf_13_wb_clk_i _01721_ _00389_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12586__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__A _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12793_ net378 _06432_ _07041_ _07316_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_194_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14532_ net1134 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11744_ net257 net2496 net596 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09671__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14463_ net1115 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XANTENNA__13204__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ _04865_ _05985_ _06531_ _07160_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16202_ clknet_leaf_37_wb_clk_i _02342_ _01010_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13414_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09959__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10626_ _06128_ _06142_ _04490_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a21oi_4
X_14394_ net1087 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10569__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output191_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16133_ clknet_leaf_28_wb_clk_i _02273_ _00941_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13345_ team_02_WB.instance_to_wrap.ramload\[7\] net1015 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[7\] sky130_fd_sc_hd__and2_1
X_10557_ _06072_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16064_ clknet_leaf_17_wb_clk_i _02204_ _00872_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13276_ net1610 net984 net966 _02987_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__a22o_1
X_10488_ _05649_ _06004_ _05624_ _05646_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11518__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15015_ net1146 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
X_12227_ net1926 net309 net613 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ net284 net1987 net462 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
X_11109_ net837 _06596_ _06617_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__o21bai_4
XPHY_EDGE_ROW_16_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12089_ net2272 net273 net583 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
XANTENNA__10789__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15917_ clknet_leaf_49_wb_clk_i _02057_ _00725_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ clknet_leaf_10_wb_clk_i _01988_ _00656_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire505_A _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12496__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15779_ clknet_leaf_10_wb_clk_i _01919_ _00587_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_08320_ _04032_ _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__nand2_1
XANTENNA__10257__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08251_ _03945_ _03957_ _03960_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10009__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11206__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08182_ _03888_ _03893_ _03862_ _03878_ _03887_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_131_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09414__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput210 net210 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput221 net221 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_11_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12182__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout487_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _03687_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__or2_1
X_09705_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\] net714 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\]
+ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ _03588_ _03598_ _03595_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09636_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\] net829 net821 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\]
+ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11307__C net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_143_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] net742 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ _04207_ net1600 net849 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_43_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09498_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\] net738 _05011_ _05013_
+ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10799__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09653__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08449_ _04153_ _03321_ net1006 net1622 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ net1695 net324 net637 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XANTENNA__09405__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ net517 _05419_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ net973 _06206_ _06885_ _06889_ _06837_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a311o_1
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13130_ _07375_ _07376_ _07415_ net976 vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a31o_1
X_10342_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] net749 net713 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ team_02_WB.instance_to_wrap.top.pc\[25\] _07349_ _02837_ _02841_ vssd1 vssd1
+ vccd1 vccd1 _01506_ sky130_fd_sc_hd__o22a_1
X_10273_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\] _04530_ net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_52_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12012_ net237 net1956 net474 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XANTENNA__08916__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__Y _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout470 net473 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_6
XFILLER_0_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout481 _07204_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_4
X_16751_ net1295 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xfanout492 _07196_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_6
X_13963_ net1244 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
X_15702_ clknet_leaf_50_wb_clk_i _01842_ _00510_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12914_ _04802_ _06150_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__o21bai_1
X_16682_ clknet_leaf_65_wb_clk_i _02799_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13894_ net1167 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XFILLER_0_186_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09892__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ clknet_leaf_128_wb_clk_i _01773_ _00441_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12845_ _05016_ _06184_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_61_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10239__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ _06825_ _06854_ _06876_ _06925_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__and4_1
X_15564_ clknet_leaf_124_wb_clk_i _01704_ _00372_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ net1079 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ net325 net2179 net601 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08852__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15495_ clknet_leaf_38_wb_clk_i _01635_ _00303_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11451__A2 _06942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ _05830_ _05908_ _05907_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__a21oi_1
X_14446_ net1073 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_211_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ net550 _04491_ _04494_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09197__Y _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ net1221 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
X_11589_ _05910_ net663 _06113_ _05783_ _07077_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold907 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16116_ clknet_leaf_3_wb_clk_i _02256_ _00924_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13328_ net1586 _03010_ _03012_ _03292_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[1\]
+ sky130_fd_sc_hd__a22o_1
Xhold918 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_70_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold929 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16047_ clknet_leaf_41_wb_clk_i _02187_ _00855_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13259_ _02964_ _02976_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07820_ _03541_ _03542_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10190__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _03471_ _03472_ _03467_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a21o_1
XANTENNA__10312__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13904__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07682_ _03393_ _03394_ _03369_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__a2111o_1
X_09421_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] net822 net818 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\]
+ _04931_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\] net740 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09096__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09635__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08303_ _04000_ _04007_ _04016_ _03992_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a31o_2
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09283_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] net779 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a221o_1
XANTENNA__08843__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ _03897_ _03922_ _03923_ _03913_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ _03880_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout402_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08096_ _03815_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand2_2
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload91 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_100_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09564__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _04295_ net945 _04507_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__and3_4
XANTENNA__10181__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ _03632_ _03634_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13236__D _04346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13814__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _06471_ _06472_ net415 vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09619_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] net738 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__a221o_1
X_10891_ net409 _06404_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ net2087 net336 net553 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__mux2_1
XANTENNA__10876__C _06080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11334__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input102_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09626__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ net319 net2359 net443 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08834__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11512_ net794 _07001_ _07002_ net654 _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__o221a_1
X_14300_ net1193 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
X_15280_ clknet_leaf_68_wb_clk_i _01424_ _00093_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ net298 net2448 net558 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ net1185 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11443_ _06896_ _06938_ net368 vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11197__A1 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14162_ net1177 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
X_11374_ net423 _06406_ _06872_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10944__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13113_ net229 _02884_ _06811_ net232 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_189_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10325_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\] net870 _05841_ vssd1
+ vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a21o_1
X_14093_ net1120 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
X_13044_ _07356_ _07357_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__nand2b_1
X_10256_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] net743 net739 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22o_1
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1221 net1222 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
Xfanout1232 net1236 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_4
XANTENNA__12104__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] net888 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a22o_1
Xfanout1243 net1264 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_4
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__buf_2
Xfanout1265 net38 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
X_14995_ net1154 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XANTENNA__11943__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16734_ net1362 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
X_13946_ net1240 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09865__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16665_ clknet_leaf_70_wb_clk_i _02784_ _01407_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13877_ net1263 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08096__Y _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15616_ clknet_leaf_109_wb_clk_i _01756_ _00424_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09078__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ team_02_WB.instance_to_wrap.top.i_ready team_02_WB.instance_to_wrap.top.testpc.en_latched
+ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__and2b_1
XFILLER_0_186_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16596_ clknet_leaf_90_wb_clk_i _02715_ _01389_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09617__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15547_ clknet_leaf_33_wb_clk_i _01687_ _00355_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08825__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ _04610_ _04653_ _04735_ _04949_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__or4_1
XANTENNA__14555__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15478_ clknet_leaf_49_wb_clk_i _01618_ _00286_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14429_ net1207 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold704 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold726 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold748 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] net676 _05483_ _05486_
+ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] net1009 _04232_ _04442_ vssd1
+ vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08852_ net142 net1042 net1034 net1392 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XANTENNA__12014__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10163__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _03481_ _03494_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nor2_1
XANTENNA_wire625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A1_N net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08783_ _04296_ _04358_ _04363_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09305__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ _03419_ _03444_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__o21a_2
XFILLER_0_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09856__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07665_ _03356_ _03357_ _03361_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout352_A _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09404_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] net779 _04917_ _04918_
+ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1094_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09069__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07596_ net1010 _03317_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nand2_2
XFILLER_0_153_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\] net810 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\]
+ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__a221o_1
XANTENNA__12612__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12684__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14465__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09266_ _04777_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08217_ _03900_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13168__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09197_ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08148_ _03863_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__nor2_1
XANTENNA__09241__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__X _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08079_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03796_ _03797_ _03798_ vssd1
+ vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__12713__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10110_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] _04326_ net650 _05626_
+ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a22oi_4
X_11090_ _05127_ _06598_ _05124_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _05534_ _05556_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2_1
XANTENNA__11351__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 net176 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _02574_ vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_02_WB.instance_to_wrap.top.a1.data\[5\] vssd1 vssd1 vccd1 vccd1 net1404
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_02_WB.instance_to_wrap.ramstore\[19\] vssd1 vssd1 vccd1 vccd1 net1415
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] vssd1 vssd1
+ vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 team_02_WB.instance_to_wrap.top.a1.data\[0\] vssd1 vssd1 vccd1 vccd1 net1437
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13800_ net1426 _03284_ _03286_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__a21oi_1
Xhold86 team_02_WB.START_ADDR_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13544__A team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold97 net164 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14780_ net1200 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
X_11992_ net310 net1828 net478 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XANTENNA__08638__A team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ net667 _06446_ _06455_ _06456_ _06428_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_202_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] _03240_ vssd1 vssd1 vccd1
+ vccd1 _03241_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08992__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16450_ clknet_leaf_62_wb_clk_i net1454 _01258_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
X_10874_ net392 _06074_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__or2_1
X_13662_ net1365 _04100_ net851 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15401_ clknet_leaf_113_wb_clk_i _01541_ _00209_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12613_ net1671 net266 net554 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__mux2_1
XANTENNA__11406__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12594__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13593_ team_02_WB.instance_to_wrap.top.a1.row2\[1\] _03126_ _03023_ vssd1 vssd1
+ vccd1 vccd1 _03147_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16381_ clknet_leaf_87_wb_clk_i _02516_ _01189_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08807__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15332_ clknet_leaf_62_wb_clk_i _01475_ _00145_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12544_ net255 net1837 net445 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15263_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[22\]
+ _00076_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_12475_ net242 net1959 net558 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
X_14214_ net1212 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
X_11426_ net414 _06483_ net423 vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09232__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 team_02_WB.instance_to_wrap.ramload\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ net1247 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08660__X _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_54_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14145_ net1261 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XANTENNA__11938__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11357_ net836 _06844_ _06856_ _06842_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10308_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\] net745 _05824_ vssd1
+ vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a21o_1
X_14076_ net1201 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
X_11288_ net606 _06783_ _06790_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_169_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10475__A_N net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _07444_ _07445_ _07446_ _07537_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__a22o_1
X_10239_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] net928 net920 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ _05755_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10145__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1040 net1046 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1062 team_02_WB.instance_to_wrap.top.a1.instruction\[5\] vssd1 vssd1 vccd1
+ vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
Xfanout1095 net1100 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_4
XFILLER_0_206_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09299__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14978_ net1154 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_109_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16717_ net1276 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
X_13929_ net1233 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16648_ clknet_leaf_92_wb_clk_i _02767_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16579_ clknet_leaf_91_wb_clk_i _02698_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\] net832 net828 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\]
+ _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09471__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09051_ net546 _04565_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03723_ _03724_ vssd1 vssd1
+ vccd1 vccd1 _03725_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold501 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09223__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10908__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold512 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold534 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13629__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold556 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\] net770 net742 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ net1047 _04187_ _04199_ net1009 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_51_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1048_A team_02_WB.instance_to_wrap.ramload\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09884_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] net812 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a22o_1
XANTENNA__10136__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1107_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1201 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1
+ net2563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ net1449 net1043 net1035 team_02_WB.instance_to_wrap.ramstore\[29\] vssd1
+ vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
Xhold1223 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10687__A3 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1234 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12679__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout567_A _07218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] net737 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a22o_1
Xhold1267 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ _03438_ _03439_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__or2_1
X_08697_ net1001 net848 vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__and2_2
XFILLER_0_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout734_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ _03342_ _03360_ _03339_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout901_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ net2561 net187 _00017_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1264_X net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12708__A _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10941__A2_N net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] net731 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10590_ _05809_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__or2_1
XANTENNA__08193__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09249_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\] _04765_ vssd1 vssd1 vccd1
+ vccd1 _04766_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14923__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13546__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12260_ net311 net1984 net575 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09214__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ _06605_ _06715_ net399 vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11758__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12191_ net285 net2063 net576 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11142_ _06178_ _06228_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__nor2_1
XANTENNA__13313__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _06104_ _06122_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__nor2_2
X_15950_ clknet_leaf_47_wb_clk_i _02090_ _00758_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10127__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\] net916 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a22o_1
X_14901_ net1200 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ clknet_leaf_116_wb_clk_i _02021_ _00689_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14832_ net1225 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XANTENNA__13077__B2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_101_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14763_ net1152 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XANTENNA__15262__Q team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ net643 _07203_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16502_ clknet_leaf_127_wb_clk_i _02636_ _01309_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_13714_ net1139 _03230_ _03231_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__nor3_1
X_10926_ _06334_ _06337_ net369 vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14694_ net1204 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16433_ clknet_leaf_44_wb_clk_i net1384 _01241_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ net2613 net245 net639 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
X_13645_ net1564 net963 _03192_ net1068 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12177__X _07214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16364_ clknet_leaf_126_wb_clk_i _02504_ _01172_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ net517 net402 vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13576_ team_02_WB.instance_to_wrap.top.a1.row1\[120\] _03116_ _03121_ team_02_WB.instance_to_wrap.top.a1.row1\[112\]
+ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10063__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ clknet_leaf_43_wb_clk_i _01458_ _00128_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10063__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ net312 net2279 net447 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
X_16295_ clknet_leaf_38_wb_clk_i _02435_ _01103_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_15246_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[5\]
+ _00059_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09205__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net311 net1812 net451 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ net836 _06895_ _06902_ _06117_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__o221a_1
X_15177_ net1145 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12389_ net286 net2034 net459 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10366__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14128_ net1232 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14059_ net1137 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XANTENNA__10118__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire535_A _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12499__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08620_ net75 net1557 net956 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10601__A _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08551_ _04208_ _04209_ net651 net792 net1596 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a32o_1
XANTENNA__11618__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12815__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ _00017_ _04170_ _04176_ _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09103_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\] net697 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout315_A _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09034_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] net912 _04530_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ _04549_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold320 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11554__A1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11554__B2 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold353 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_8
Xhold386 team_02_WB.instance_to_wrap.top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1 net1748
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15368__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold397 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net1759 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 _04522_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08970__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\] net812 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\]
+ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a221o_1
Xfanout822 _04514_ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_8
Xfanout833 _04506_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_2
Xfanout844 _04400_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_8
Xfanout855 _04550_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_8
Xfanout866 net869 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_181_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 _04539_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] net765 net753 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\]
+ _05383_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a221o_1
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_4
XFILLER_0_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1020 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 _04526_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_2
Xhold1042 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] vssd1
+ vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12202__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ net1519 net1040 net993 team_02_WB.instance_to_wrap.ramaddr\[13\] vssd1 vssd1
+ vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09798_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] net896 net943 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a22o_1
Xhold1064 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08749_ _04296_ _04359_ _04370_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14918__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ net321 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\] net596 vssd1
+ vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__mux2_1
XANTENNA__09683__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _06181_ _06227_ _06182_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _05738_ _05916_ _07141_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11342__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13430_ _03038_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__inv_2
X_10642_ _04268_ _06155_ _06157_ _04311_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__o22a_1
XANTENNA__09435__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13231__B2 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ net2514 net1016 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[23\]
+ sky130_fd_sc_hd__and2_1
X_10573_ _05187_ net386 _06089_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14653__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15100_ net1105 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
X_12312_ net238 net1710 net564 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__mux2_1
X_16080_ clknet_leaf_23_wb_clk_i _02220_ _00888_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13292_ net1614 net984 net966 _02995_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__a22o_1
XANTENNA_input78_A wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12243_ _04291_ net643 _07188_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__or3_1
X_15031_ net1244 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XANTENNA__10348__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12174_ net363 net1807 net462 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16293__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net409 _06347_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__nand2_1
XANTENNA__09753__Y _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13298__B2 _02998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ _05950_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nor2_1
X_15933_ clknet_leaf_13_wb_clk_i _02073_ _00741_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10007_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] net696 _05521_ _05523_
+ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a211o_1
XANTENNA__11517__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_199_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ clknet_leaf_121_wb_clk_i _02004_ _00672_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12112__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ net1116 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15795_ clknet_leaf_59_wb_clk_i _01935_ _00603_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11951__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13291__X _02995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ net1087 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09674__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__A1 team_02_WB.START_ADDR_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11958_ net309 net2521 net585 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10909_ _06419_ _06423_ net605 _06416_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__o211a_4
XFILLER_0_74_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14677_ net1242 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
X_11889_ net300 net2028 net488 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16416_ clknet_leaf_99_wb_clk_i _02551_ _01224_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_15_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13628_ team_02_WB.instance_to_wrap.top.a1.row1\[60\] _03117_ _03160_ team_02_WB.instance_to_wrap.top.a1.row1\[108\]
+ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__a221o_1
XANTENNA__09426__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16347_ clknet_leaf_32_wb_clk_i _02487_ _01155_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13559_ net1052 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] vssd1 vssd1 vccd1
+ vccd1 _03114_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ clknet_leaf_22_wb_clk_i _02418_ _01086_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15510__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15229_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[20\]
+ _00042_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11536__A1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07982_ _03677_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__or2_1
XANTENNA__13289__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\] net799 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12022__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\] net783 net759 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a22o_1
X_08603_ net93 net1414 net957 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
X_09583_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\] net698 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16016__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ _04219_ net1669 net849 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09665__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11472__B1 _06965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] _04158_ _04160_ vssd1 vssd1
+ vccd1 vccd1 _04166_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1174_A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09417__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04070_ vssd1 vssd1 vccd1
+ vccd1 _04105_ sky130_fd_sc_hd__xor2_2
XFILLER_0_135_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire508 _05578_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_2
Xwire519 _05313_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13285__A1_N _06782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09838__Y _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08471__A team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout899_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _04510_ _04516_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__nor2_4
XFILLER_0_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold150 team_02_WB.START_ADDR_VAL_REG\[25\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold161 team_02_WB.START_ADDR_VAL_REG\[26\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_02_WB.START_ADDR_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_02_WB.instance_to_wrap.ramstore\[29\] vssd1 vssd1 vccd1 vccd1 net1545
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 team_02_WB.instance_to_wrap.top.a1.row1\[11\] vssd1 vssd1 vccd1 vccd1 net1556
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13817__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout641 _04453_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_6
XFILLER_0_186_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09919_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\] net733 net677 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__a22o_1
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 _06111_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net676 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_8
Xfanout685 _04399_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_4
Xfanout696 _04394_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ team_02_WB.instance_to_wrap.top.pc\[28\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _07450_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_161_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ net515 _05444_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__or2_1
X_14600_ net1112 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
X_11812_ net265 net2490 net590 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15580_ clknet_leaf_20_wb_clk_i _01720_ _00388_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12792_ _06054_ _06296_ net384 vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11463__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ net1133 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XANTENNA__09120__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11743_ net248 net2412 net597 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09408__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14462_ net1191 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
X_11674_ _06373_ _07158_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ clknet_leaf_111_wb_clk_i _02341_ _01009_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11215__B1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] net995 vssd1 vssd1 vccd1
+ vccd1 _06142_ sky130_fd_sc_hd__nand2_1
X_14393_ net1095 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16132_ clknet_leaf_36_wb_clk_i _02272_ _00940_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09477__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10556_ _04802_ net405 vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__nor2_1
XANTENNA__08092__C1 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ net2249 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[6\]
+ sky130_fd_sc_hd__and2_1
X_16063_ clknet_leaf_58_wb_clk_i _02203_ _00871_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10487_ _05913_ _06003_ _05914_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__a21o_1
XANTENNA__12107__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13275_ _06648_ _02959_ team_02_WB.instance_to_wrap.top.pc\[22\] net1055 vssd1 vssd1
+ vccd1 vccd1 _02987_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_121_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11518__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15014_ net1162 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XANTENNA__09187__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ net2106 net303 net615 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_184_Right_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11946__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ net272 net2112 net464 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
X_11108_ net671 _06603_ _06609_ _06104_ _06616_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__a221o_1
X_12088_ net2242 net290 net581 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
X_11039_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__inv_2
X_15916_ clknet_leaf_2_wb_clk_i _02056_ _00724_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10151__A team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15847_ clknet_leaf_38_wb_clk_i _01987_ _00655_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15778_ clknet_leaf_116_wb_clk_i _01918_ _00586_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08556__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09111__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__X _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ net1222 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08250_ _03956_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_31_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ _03886_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_41_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08622__A1 team_02_WB.START_ADDR_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12017__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput211 net211 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput222 net222 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_140_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11856__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13196__X _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10193__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__X _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07635__A team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07965_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03670_ _03672_ vssd1 vssd1
+ vccd1 vccd1 _03688_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09704_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\] net742 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07896_ net316 _03597_ _03588_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a21o_1
XANTENNA__09886__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09350__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09635_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] net817 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a22o_1
XANTENNA__12687__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09566_ _05082_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__inv_2
XANTENNA__09638__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09102__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ net1048 _04205_ _04206_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\] net786 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout814_A _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _04149_ _04150_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08753__X _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _04084_ _04085_ _04081_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07962__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10410_ _05468_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11390_ _06200_ net652 _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] _06888_
+ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__a221o_1
XANTENNA__09810__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\] net769 net745 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14931__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09169__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ _04280_ _02839_ _02840_ net230 net1026 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a221o_1
X_10272_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] net824 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ net244 net2401 net476 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11619__X _07107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10184__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 _07220_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_6
Xfanout471 net473 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_8
X_16750_ net1294 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
Xfanout482 _07200_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_6
Xfanout493 _07196_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_4
X_13962_ net1244 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
X_15701_ clknet_leaf_31_wb_clk_i _01841_ _00509_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09341__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12913_ _04842_ _06172_ _07432_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__a21oi_1
X_16681_ clknet_leaf_65_wb_clk_i _02798_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12597__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ net1166 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ clknet_leaf_23_wb_clk_i _01772_ _00440_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12844_ _04971_ _06180_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15563_ clknet_leaf_15_wb_clk_i _01703_ _00371_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12775_ _06360_ _06452_ _07297_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__and4_1
XFILLER_0_185_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15270__Q team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ net1184 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
X_11726_ net323 net1760 net600 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15494_ clknet_leaf_10_wb_clk_i _01634_ _00302_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14445_ net1121 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
X_11657_ _05832_ _05910_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14376_ net1104 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XANTENNA__09801__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _05909_ net657 vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16115_ clknet_leaf_56_wb_clk_i _02255_ _00923_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold908 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ _00009_ team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] vssd1 vssd1 vccd1
+ vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] sky130_fd_sc_hd__or2_1
Xmax_cap616 net617 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10539_ _05489_ net403 vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__or2_1
Xhold919 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net2281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14841__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16046_ clknet_leaf_46_wb_clk_i _02186_ _00854_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13258_ _06458_ _02963_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__and2_1
X_12209_ net347 net2499 net576 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13189_ _04280_ _07395_ _02945_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a31o_1
XFILLER_0_193_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07750_ _03471_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__nand2_1
XANTENNA__09868__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ _03393_ _03394_ _03369_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09420_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\] net814 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12300__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09351_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\] net788 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a22o_1
X_08302_ _04000_ _04007_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09282_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\] net751 net739 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08233_ _03913_ _03927_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09399__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ _03840_ net227 _03847_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08095_ _03782_ _03786_ _03811_ _03785_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout1137_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_2
Xclkload81 clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_8
XFILLER_0_100_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload92 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload92/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout597_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__A net2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11439__X _06936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10166__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09571__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10062__Y _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _04297_ net944 _04503_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_145_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10602__A2_N _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ _03631_ _03634_ _03637_ _03622_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__a31o_1
XANTENNA__09859__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09323__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07879_ _03571_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09618_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\] net690 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__a22o_1
X_10890_ _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09549_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\] net814 net810 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ net312 net1889 net442 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ net665 _06053_ net378 _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_199_Left_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08771__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12491_ net310 net2064 net557 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ net1107 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
X_11442_ _06301_ _06304_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ net375 _06665_ _06871_ net380 vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__o22a_1
X_14161_ net1232 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09177__D _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input60_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\] net910 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a22o_1
X_13112_ _07516_ _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_189_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14092_ net1216 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13043_ team_02_WB.instance_to_wrap.top.pc\[28\] _07349_ _02822_ _02826_ vssd1 vssd1
+ vccd1 vccd1 _01509_ sky130_fd_sc_hd__o22a_1
X_10255_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] net715 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a221o_1
XANTENNA__10157__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1211 net1237 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_2
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_4
X_10186_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] net807 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__a221o_1
Xfanout1233 net1235 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
XANTENNA__15265__Q team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1244 net1249 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_208_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1255 net1264 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_2
X_14994_ net1133 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09314__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16733_ net1361 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
X_13945_ net1255 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11525__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12120__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ clknet_leaf_93_wb_clk_i _02783_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13876_ net1250 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
XFILLER_0_186_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15615_ clknet_leaf_59_wb_clk_i _01755_ _00423_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11409__B1 _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ team_02_WB.instance_to_wrap.top.a1.state\[0\] _07343_ _07345_ _07347_ vssd1
+ vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__o22a_1
X_16595_ clknet_leaf_97_wb_clk_i _02714_ _01388_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14836__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ clknet_leaf_52_wb_clk_i _01686_ _00354_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12758_ _05648_ _05915_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11709_ net251 net1890 net602 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15477_ clknet_leaf_49_wb_clk_i _01617_ _00285_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12689_ net310 net1686 net431 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14428_ net1199 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold705 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ net1185 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XANTENNA__14571__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_203_Left_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold716 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold749 team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] vssd1 vssd1 vccd1 vccd1
+ net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12803__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] net958 _04212_ _04173_ vssd1
+ vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o211a_1
X_16029_ clknet_leaf_12_wb_clk_i _02169_ _00837_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09002__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10148__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11896__A0 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ net143 net1043 net1035 net1398 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
XANTENNA__09553__A2 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11419__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13915__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _03512_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__and2_1
X_08782_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] net753 net709 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\]
+ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__A2 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07733_ _03413_ _03416_ _03445_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a31o_1
XANTENNA__11112__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12030__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07664_ _03384_ _03385_ _03351_ _03383_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and4b_1
XANTENNA__10320__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09403_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\] net727 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\]
+ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07595_ net1010 _03317_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout345_A _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1087_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\] net925 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09265_ net536 _04775_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__nand2_1
XANTENNA__10338__X _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _03884_ _03899_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09196_ _04702_ _04707_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__nor3_4
XFILLER_0_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11179__A2 _06679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08147_ _03829_ net227 _03835_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__C1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09792__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ _03797_ _03798_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout881_A _04538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15744__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10040_ _05534_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 team_02_WB.instance_to_wrap.top.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 net1372
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_02_WB.instance_to_wrap.ramstore\[6\] vssd1 vssd1 vccd1 vccd1 net1383
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 team_02_WB.instance_to_wrap.ramstore\[5\] vssd1 vssd1 vccd1 vccd1 net1394
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net182 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _02581_ vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold65 net130 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net179 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net160 vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11616__Y _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13544__B _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 _02565_ vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11991_ net300 net2589 net479 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ _03240_ net951 _03239_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__and3b_1
X_10942_ _04693_ net661 _06453_ net795 vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_67_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13661_ net1368 _04111_ net851 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10873_ _06382_ _06387_ net412 vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15400_ clknet_leaf_25_wb_clk_i _01540_ _00208_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12612_ net2304 net260 net552 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__mux2_1
X_16380_ clknet_leaf_84_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[4\] _01188_
+ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__dfrtp_1
X_13592_ team_02_WB.instance_to_wrap.top.a1.row1\[57\] _03117_ _03119_ team_02_WB.instance_to_wrap.top.a1.row1\[1\]
+ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_80_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ clknet_leaf_62_wb_clk_i _01474_ _00144_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11351__Y _06851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12543_ net238 net2447 net442 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
X_15262_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[21\]
+ _00075_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10090__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12474_ _04292_ _04452_ _07201_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__or3_4
X_14213_ net1113 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
X_11425_ net376 _06716_ _06921_ net382 vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15193_ net1247 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_14144_ net1104 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XANTENNA__09783__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ net666 _06845_ _06852_ _06855_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_111_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] net717 net701 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a22o_1
X_14075_ net1087 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XANTENNA__12115__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ net973 _06784_ _06789_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_169_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09535__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13026_ _07444_ _07445_ _07446_ _07537_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__nand4_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\] net884 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_206_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_206_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11954__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1041 net1046 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1052 team_02_WB.instance_to_wrap.top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1
+ net1052 sky130_fd_sc_hd__dlymetal6s2s_1
X_10169_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\] net876 _05675_ _05685_
+ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a211o_1
Xfanout1063 team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1 vccd1
+ vccd1 net1063 sky130_fd_sc_hd__buf_2
Xfanout1074 net1101 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_4
XFILLER_0_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1100 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__buf_4
X_14977_ net1154 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_109_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13928_ net1228 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
X_16716_ net1275 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XANTENNA__10302__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16647_ clknet_leaf_92_wb_clk_i _02766_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13859_ net1151 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16578_ clknet_leaf_91_wb_clk_i _00004_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09012__X _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15529_ clknet_leaf_110_wb_clk_i _01669_ _00337_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ net546 _04565_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10081__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__X _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ _03305_ net256 _03689_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15767__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10369__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold513 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11030__A1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold535 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10605__Y _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] vssd1 vssd1
+ vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12025__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__inv_2
Xhold579 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09526__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08903_ team_02_WB.instance_to_wrap.top.edg2.flip2 _04179_ _04182_ team_02_WB.instance_to_wrap.top.edg2.flip1
+ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_148_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09883_ _05384_ _05390_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_5_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11864__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_148_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08834_ net162 net1042 net1034 net1386 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
Xhold1213 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1224 team_02_WB.instance_to_wrap.top.d_ready vssd1 vssd1 vccd1 vccd1 net2586
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07643__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1246 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13364__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ net846 _04363_ _04364_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout462_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1268 team_02_WB.instance_to_wrap.top.a1.row1\[60\] vssd1 vssd1 vccd1 vccd1 net2630
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07716_ _03403_ net425 _03408_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ _04323_ _04324_ _04307_ _04322_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_196_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07647_ _03343_ _03360_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nor2_2
XANTENNA__12695__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15297__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__nor2_1
XFILLER_0_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09317_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] net675 _04824_ _04827_
+ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09248_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a22o_1
XANTENNA__10072__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09179_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\] net727 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a22o_1
XANTENNA__16692__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _06662_ _06714_ net370 vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__mux2_1
X_12190_ net273 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] net579 vssd1
+ vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_1
XANTENNA__09765__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ net954 _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nand2_1
XANTENNA__10244__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11072_ _04864_ net659 _06122_ _06357_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__a22o_1
XANTENNA__09517__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput100 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
X_10023_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] net929 net885 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a221o_1
XANTENNA__11774__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14900_ net1153 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
X_15880_ clknet_leaf_20_wb_clk_i _02020_ _00688_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14831_ net1219 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14762_ net1177 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11974_ _07188_ _07201_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_201_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09150__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ clknet_leaf_0_wb_clk_i _02635_ _01308_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13713_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\]
+ _03227_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__and3_1
X_10925_ _06309_ _06331_ net369 vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_127_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14693_ net1172 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XANTENNA__08655__Y _04284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16432_ clknet_leaf_61_wb_clk_i net1395 _01240_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
X_13644_ _03023_ _03185_ _03189_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or4_1
X_10856_ net946 _06365_ _06371_ net604 vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__o211a_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ clknet_leaf_14_wb_clk_i _02503_ _01171_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13575_ team_02_WB.instance_to_wrap.top.a1.row2\[40\] _03123_ _03125_ team_02_WB.instance_to_wrap.top.a1.row2\[32\]
+ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10419__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ _06299_ _06302_ net367 vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__mux2_1
X_15314_ clknet_leaf_44_wb_clk_i _01457_ _00127_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12526_ net305 net2182 net449 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
XANTENNA__10063__A2 _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16294_ clknet_leaf_6_wb_clk_i _02434_ _01102_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11949__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13289__X _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15245_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[4\]
+ _00058_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12457_ net301 net1778 net452 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15010__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _06037_ _06903_ _06905_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09756__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15176_ net1143 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_136_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12388_ net272 net2476 net460 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14127_ net1224 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
X_11339_ net948 _06830_ _06839_ net607 vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__o211a_4
XANTENNA__09508__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14058_ net1118 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13009_ team_02_WB.instance_to_wrap.top.pc\[23\] _06177_ _07528_ vssd1 vssd1 vccd1
+ vccd1 _07529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_207_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09007__X _04524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08550_ _04205_ _04206_ _04224_ net793 net1659 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_145_Left_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09141__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08481_ team_02_WB.instance_to_wrap.top.a1.state\[0\] _04168_ vssd1 vssd1 vccd1 vccd1
+ _04180_ sky130_fd_sc_hd__nand2_2
XFILLER_0_76_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12809__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09102_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] net769 net701 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10054__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_198_Right_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09033_ net945 _04528_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__nor2_4
XANTENNA__11859__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_Left_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold310 team_02_WB.instance_to_wrap.top.a1.row1\[114\] vssd1 vssd1 vccd1 vccd1 net1672
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09747__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1158_A team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold365 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold376 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1217_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 team_02_WB.instance_to_wrap.top.a1.row2\[12\] vssd1 vssd1 vccd1 vccd1 net1749
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _04535_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_4
X_09935_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] net926 net922 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a22o_1
Xfanout812 net813 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
Xfanout823 _04514_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 _04506_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout677_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__X _06943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 _04400_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13375__A net2352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13700__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 _04550_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
X_09866_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] net777 net717 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a22o_1
Xfanout867 net869 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_181_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 _04538_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1010 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _04536_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_8
Xhold1032 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net1498 net1041 net991 team_02_WB.instance_to_wrap.ramaddr\[14\] vssd1 vssd1
+ vccd1 vccd1 _02608_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_163_Left_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1043 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ net519 vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__inv_2
XANTENNA__15363__Q team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1054 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _04302_ net847 _04365_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__and3_1
Xhold1098 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08756__X _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_X clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ net1063 _04266_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__and2_1
XANTENNA__15932__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10710_ team_02_WB.instance_to_wrap.top.pc\[20\] _06184_ _06226_ vssd1 vssd1 vccd1
+ vccd1 _06227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10293__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11690_ _07140_ _07143_ _07161_ _07175_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08635__C team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10641_ _04272_ _04277_ _04276_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13231__A2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ net2520 net1016 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[22\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_146_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10572_ net524 net386 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_172_Left_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09986__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ net244 net2058 net565 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__mux2_1
XANTENNA__11769__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ _06857_ _02959_ team_02_WB.instance_to_wrap.top.pc\[14\] net1056 vssd1 vssd1
+ vccd1 vccd1 _02995_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08651__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09199__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15030_ net1250 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
X_12242_ net1934 net349 net612 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__mux2_1
XANTENNA__09738__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08946__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12173_ net354 net2575 net464 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11124_ net409 _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_166_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13298__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__X _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11055_ _04865_ _05949_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__nor2_1
X_15932_ clknet_leaf_17_wb_clk_i _02072_ _00740_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_181_Left_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09371__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\] net844 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\]
+ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__a221o_1
XANTENNA_input26_X net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09910__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15863_ clknet_leaf_120_wb_clk_i _02003_ _00671_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_199_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14814_ net1188 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
X_15794_ clknet_leaf_56_wb_clk_i _01934_ _00602_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14745_ net1091 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
X_11957_ net301 net1887 net586 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10284__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11481__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ net999 _06422_ _06420_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14676_ net1238 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
X_11888_ net294 net1862 net487 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
X_16415_ clknet_leaf_99_wb_clk_i _02550_ _01223_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[22\]
+ sky130_fd_sc_hd__dfrtp_2
X_13627_ team_02_WB.instance_to_wrap.top.a1.row1\[12\] _03109_ _03114_ _03177_ vssd1
+ vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a31o_1
X_10839_ net545 net424 vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_15_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14844__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16346_ clknet_leaf_50_wb_clk_i _02486_ _01154_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13558_ net1051 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] vssd1 vssd1 vccd1
+ vccd1 _03113_ sky130_fd_sc_hd__nor2_2
XANTENNA__09977__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ net244 net2080 net448 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__mux2_1
XANTENNA__10583__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16277_ clknet_leaf_22_wb_clk_i _02417_ _01085_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13489_ team_02_WB.START_ADDR_VAL_REG\[29\] _04260_ vssd1 vssd1 vccd1 vccd1 net213
+ sky130_fd_sc_hd__and2_1
XFILLER_0_120_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15228_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[19\]
+ _00041_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09729__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15159_ net1144 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XANTENNA_max_cap528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07981_ _03698_ net256 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_130_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13289__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] net919 net805 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\]
+ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a221o_1
XANTENNA__10612__A team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12303__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net525 _05165_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08602_ net95 net1539 net955 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
X_09582_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] net765 net729 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08533_ _04171_ _04217_ _04218_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout258_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11472__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ net1560 net1006 net981 _04165_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
XANTENNA__11472__B2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _04095_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14754__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1167_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09968__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09016_ net945 _04505_ _04509_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10065__Y _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold140 _02564_ vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold151 team_02_WB.START_ADDR_VAL_REG\[21\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 team_02_WB.START_ADDR_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 team_02_WB.START_ADDR_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold184 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_02_WB.START_ADDR_VAL_REG\[12\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\] net769 net717 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a22o_1
XANTENNA__12488__A0 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout642 _04453_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_2
XANTENNA__12213__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 _06247_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10522__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 _06111_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
XANTENNA__13205__A2_N net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout686 _04399_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout697 _04391_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_8
X_09849_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\] net825 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a22o_1
XANTENNA__11337__B _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ net518 _07378_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_161_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08927__A team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11811_ net257 net2229 net588 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791_ _06612_ _06641_ _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__and3_1
XFILLER_0_201_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14530_ net1152 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11742_ net254 net1902 net599 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14461_ net1203 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
X_11673_ _04783_ _06467_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16200_ clknet_leaf_20_wb_clk_i _02340_ _01008_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13412_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _03024_
+ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input90_A wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09959__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ team_02_WB.instance_to_wrap.top.pc\[28\] _06139_ vssd1 vssd1 vccd1 vccd1
+ _06141_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14392_ net1189 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
X_16131_ clknet_leaf_25_wb_clk_i _02271_ _00939_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13343_ team_02_WB.instance_to_wrap.ramload\[5\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[5\] sky130_fd_sc_hd__and2_1
X_10555_ _04842_ net387 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_77_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16062_ clknet_leaf_5_wb_clk_i _02202_ _00870_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13274_ net1627 net985 net967 _02986_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net417 net501 _05738_ _06002_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o22a_1
XANTENNA__15268__Q team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15013_ net1162 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11518__A2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ net1705 net292 net612 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09592__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net288 net1994 net462 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XANTENNA__08601__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ net667 _06612_ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12123__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net1788 net276 net580 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XANTENNA__09344__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ _05809_ _06403_ _06545_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a21oi_2
X_15915_ clknet_leaf_14_wb_clk_i _02055_ _00723_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10151__B _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15846_ clknet_leaf_7_wb_clk_i _01986_ _00654_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_201_Right_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15777_ clknet_leaf_103_wb_clk_i _01917_ _00585_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12989_ _07480_ _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11454__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10257__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11454__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14728_ net1114 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14659_ net1133 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10009__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11206__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08180_ _03888_ _03893_ _03862_ _03878_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09020__X _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08083__B1 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16329_ clknet_leaf_112_wb_clk_i _02469_ _01137_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput212 net212 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XANTENNA__12706__A1 team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput223 net223 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XANTENNA__09583__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ _03670_ _03672_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1
+ vccd1 vccd1 _03687_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09335__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] net738 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__a22o_1
X_07895_ _03614_ _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14749__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] net928 net814 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\]
+ _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09565_ _05061_ _05080_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_143_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\] net979 vssd1 vssd1 vccd1
+ vccd1 _04206_ sky130_fd_sc_hd__or2_1
XANTENNA__10248__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__B2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\] net774 net757 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\]
+ _05012_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08447_ _04141_ _04146_ _04151_ _04136_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout807_A _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _04081_ _04086_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12208__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10340_ net389 vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10271_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09574__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ net242 net1899 net476 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16795__1339 vssd1 vssd1 vccd1 vccd1 _16795__1339/HI net1339 sky130_fd_sc_hd__conb_1
Xfanout450 _07222_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_6
XANTENNA__09326__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout461 _07220_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_4
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_8
X_13961_ net1167 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
Xfanout483 _07200_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_2
XANTENNA__11782__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15700_ clknet_leaf_3_wb_clk_i _01840_ _00508_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12912_ _07360_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__and2_1
X_16680_ clknet_leaf_65_wb_clk_i _02797_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13892_ net1167 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XANTENNA__11354__Y _06854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15631_ clknet_leaf_42_wb_clk_i _01771_ _00439_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _04928_ _06177_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15562_ clknet_leaf_38_wb_clk_i _01702_ _00370_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10239__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ _06482_ _06517_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__nor2_1
X_14513_ net1233 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_48_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11725_ net318 net2316 net600 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ clknet_leaf_30_wb_clk_i _01633_ _00301_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08852__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13189__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444_ net1209 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11656_ net368 _06287_ _05877_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10607_ _05962_ _06036_ _06121_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__or3_4
XFILLER_0_24_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14375_ net1174 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XANTENNA__12118__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ net378 _06470_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16114_ clknet_leaf_53_wb_clk_i _02254_ _00922_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13326_ _03292_ _03011_ _03010_ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] vssd1
+ vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] sky130_fd_sc_hd__a2bb2o_1
Xhold909 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ net509 net403 vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__nand2_1
Xmax_cap617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_2
Xmax_cap628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11957__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16045_ clknet_leaf_47_wb_clk_i _02185_ _00853_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13297__X _02998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ net1431 net983 net965 _02975_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__a22o_1
X_10469_ _05231_ _05251_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__or2_1
X_12208_ net350 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\] net576 vssd1
+ vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13188_ _07084_ net233 net230 _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10175__B2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ net356 net2416 net468 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13113__B2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07680_ _03399_ _03400_ _03402_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__a21o_1
XFILLER_0_204_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09015__X _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15829_ clknet_leaf_31_wb_clk_i _01969_ _00637_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09350_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\] net755 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09096__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08301_ _04009_ _04014_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__nor3_1
X_09281_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\] net763 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\]
+ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a221o_1
XANTENNA__08843__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ _03943_ _03944_ _03946_ _03935_ _03919_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__13222__A1_N net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08163_ _03806_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12028__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ _03801_ _03808_ _03812_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11867__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload60 clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_8
XFILLER_0_101_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload71 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload82 clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1032_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload93/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09556__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08996_ _04313_ net945 _04507_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__and3_4
XANTENNA__09308__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _03641_ _03661_ _03662_ _03663_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a41o_2
XANTENNA__09859__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12698__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__A team_02_WB.instance_to_wrap.ramload\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10800__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _03574_ _03599_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_183_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09617_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\] net706 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16694__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout924_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09548_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] net928 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a22o_1
XANTENNA__09087__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_195_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _04993_ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08834__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _05921_ net657 _05923_ net663 vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11631__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15103__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ net301 net2114 net558 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _05468_ _06009_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_22_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14942__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ net1256 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
X_11372_ _06870_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11777__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ _07468_ _07469_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nor2_1
X_10323_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] net890 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\]
+ _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14091_ net1100 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_189_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input53_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ net230 _02824_ _02825_ _04280_ net1027 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a221o_1
X_10254_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\] net687 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a22o_1
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_4
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__buf_4
Xfanout1223 net1237 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_2
X_10185_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] net822 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_208_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1245 net1249 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1256 net1262 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
XANTENNA__11106__B1 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _06657_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
X_14993_ net1135 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
Xfanout291 _06712_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11365__X _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ net1360 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__12401__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ net1255 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16663_ clknet_leaf_95_wb_clk_i _02782_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13875_ net1164 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11409__A1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15614_ clknet_leaf_4_wb_clk_i _01754_ _00422_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12826_ _07346_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__inv_2
XFILLER_0_186_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11409__B2 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09078__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16594_ clknet_leaf_89_wb_clk_i _02713_ _01387_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12757_ _05737_ _05831_ _05909_ _07128_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__or4b_1
XANTENNA__12082__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15545_ clknet_leaf_124_wb_clk_i _01685_ _00353_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10093__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11708_ net254 net1789 net602 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15476_ clknet_leaf_3_wb_clk_i _01616_ _00284_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12688_ net302 net2320 net433 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08038__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14427_ net1076 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
X_11639_ net948 _07122_ _07125_ net607 vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o211a_4
XFILLER_0_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13031__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14852__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09786__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ net1120 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XANTENNA__09250__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold717 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13468__A team_02_WB.START_ADDR_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13309_ team_02_WB.instance_to_wrap.top.pc\[5\] net1054 _07046_ net933 vssd1 vssd1
+ vccd1 vccd1 _03004_ sky130_fd_sc_hd__a22o_1
Xhold728 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ net1222 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16028_ clknet_leaf_19_wb_clk_i _02168_ _00836_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09002__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ net144 net1042 net1034 net1396 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07801_ _03519_ _03520_ _03492_ _03517_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__and4b_1
XFILLER_0_137_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08781_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\] net757 net729 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11648__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ _03423_ _03454_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__nor2_1
XANTENNA__12311__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15696__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09710__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08728__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\] net746 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09069__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ net1008 _03317_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\] net815 net912 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\]
+ _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_X clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13270__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10766__S net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16794__1338 vssd1 vssd1 vccd1 vccd1 _16794__1338/HI net1338 sky130_fd_sc_hd__conb_1
X_09264_ net536 _04776_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _03902_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09195_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] net767 _04709_ _04710_
+ _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13022__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _03833_ _03863_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09241__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13378__A team_02_WB.instance_to_wrap.ramload\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08077_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03762_ _03787_ vssd1 vssd1
+ vccd1 vccd1 _03798_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout874_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__B1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1202_X net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 _00011_ vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 _02568_ vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 _02567_ vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 team_02_WB.instance_to_wrap.top.a1.data\[1\] vssd1 vssd1 vccd1 vccd1 net1406
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net1063 net1062 _04267_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__a21o_2
XANTENNA__13089__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 team_02_WB.instance_to_wrap.ramstore\[1\] vssd1 vssd1 vccd1 vccd1 net1417
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _02625_ vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12221__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11639__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 team_02_WB.instance_to_wrap.ramaddr\[5\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 _02591_ vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net294 net2339 net480 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
Xhold99 team_02_WB.instance_to_wrap.ramaddr\[26\] vssd1 vssd1 vccd1 vccd1 net1461
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09701__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _04694_ net658 _04695_ _06111_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_203_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660_ _04125_ net851 _03197_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a21oi_1
X_10872_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ net2073 net250 net554 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13591_ team_02_WB.instance_to_wrap.top.a1.row1\[9\] _03110_ _03111_ team_02_WB.instance_to_wrap.top.a1.row1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__a22o_1
XANTENNA__08807__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08654__B team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15330_ clknet_leaf_44_wb_clk_i _01473_ _00143_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10075__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ net246 net2606 net444 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[20\]
+ _00074_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_12473_ net348 net1979 net450 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08941__Y _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14212_ net1132 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11424_ _06819_ _06920_ net396 vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__mux2_1
XANTENNA__09768__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15192_ net1141 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XANTENNA__09232__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__A team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14143_ net1108 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
X_11355_ _05295_ net664 net656 _06854_ _06846_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10306_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\] net777 net765 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a22o_1
X_14074_ net1095 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11286_ _06190_ net652 _06788_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__a21o_1
X_13025_ _06368_ net233 vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_169_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ _05747_ _05749_ _05751_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__or4_1
XANTENNA__09772__Y _05289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_2
Xfanout1031 _04430_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_2
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_2
XANTENNA__09940__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1053 team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1053 sky130_fd_sc_hd__clkbuf_4
X_10168_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\] net942 net891 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1075 net1077 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_4
Xfanout1086 net1101 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_2
XANTENNA__10440__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1100 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14976_ net1160 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
X_10099_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\] net677 _05605_ _05608_
+ _05615_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09299__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16715_ net1274 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_63_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13927_ net1244 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XANTENNA__11970__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_179_Right_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16646_ clknet_leaf_93_wb_clk_i _02765_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13858_ net1151 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12809_ net790 _07332_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nand2_1
X_16577_ clknet_leaf_92_wb_clk_i _00003_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13789_ _03278_ _03279_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15528_ clknet_leaf_24_wb_clk_i _01668_ _00336_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09471__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15459_ clknet_leaf_27_wb_clk_i _01599_ _00267_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08000_ _03689_ net256 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__nand2_1
XANTENNA__09759__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09223__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13198__A _02953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold525 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12306__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold536 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09951_ _05465_ _05466_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__nor2_2
Xhold558 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold569 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ net2 net1030 net987 net2397 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09882_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\] net725 _05391_ _05392_
+ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_51_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12830__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ net163 net1042 net1034 net1400 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a22o_1
XANTENNA__09931__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1203 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1214 team_02_WB.instance_to_wrap.top.testpc.en_latched vssd1 vssd1 vccd1 vccd1
+ net2576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] vssd1 vssd1 vccd1 vccd1
+ net2587 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout288_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] net717 _04390_ _04392_
+ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a211o_1
XANTENNA__12041__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1247 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_02_WB.instance_to_wrap.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net2631
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ _03408_ net425 _03403_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__and3b_1
XFILLER_0_79_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08695_ net1060 _03298_ _04271_ _04318_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout455_A _07221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _03363_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13380__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ team_02_WB.instance_to_wrap.top.pad.keyCode\[5\] net188 _00017_ vssd1 vssd1
+ vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\] net719 _04829_ _04830_
+ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10057__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09462__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _04757_ _04759_ _04761_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__or4_2
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1152_X net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09178_ _04693_ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09214__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout991_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08129_ _03829_ _03836_ _03837_ _03848_ _03807_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10525__A _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12216__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140_ _04470_ _06627_ _06647_ net669 _06646_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__o221a_2
XFILLER_0_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__B _05760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _04865_ _06110_ net661 _04863_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput101 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
X_10022_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] net912 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a22o_1
XANTENNA__13053__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1075 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14761_ net1222 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
X_11973_ net349 net2292 net584 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__mux2_1
XANTENNA__08489__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10296__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16500_ clknet_leaf_0_wb_clk_i _02634_ _01307_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ _06432_ _06437_ net412 vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__mux2_1
X_13712_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03227_ net1759 vssd1
+ vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__a21oi_1
X_14692_ net1098 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ clknet_leaf_44_wb_clk_i net1452 _01239_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_197_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13643_ team_02_WB.instance_to_wrap.top.a1.row1\[111\] _03160_ _03161_ _03190_ vssd1
+ vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a211o_1
XANTENNA__13234__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ net975 _06366_ _06369_ _06370_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__a211o_1
XFILLER_0_168_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10048__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16362_ clknet_leaf_39_wb_clk_i _02502_ _01170_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13574_ team_02_WB.instance_to_wrap.top.a1.row2\[8\] _03122_ _03126_ team_02_WB.instance_to_wrap.top.a1.row2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22o_1
XANTENNA__08952__X _04469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ _06300_ _06301_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__or2_1
X_15313_ clknet_leaf_45_wb_clk_i _01456_ _00126_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12525_ net296 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] net448 vssd1
+ vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__mux2_1
XANTENNA__11260__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16293_ clknet_leaf_30_wb_clk_i _02433_ _01101_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12474__X _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[3\]
+ _00057_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_12456_ net293 net2486 net451 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08604__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09205__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11407_ _05381_ _06110_ _06901_ _06104_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__a221o_1
X_15175_ net1143 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12126__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ net290 net2629 net459 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14126_ net1082 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ net973 _06212_ _06831_ _06838_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11965__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ net1228 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
X_11269_ _06714_ _06771_ net370 vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__mux2_1
X_13008_ _07457_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__and2b_1
X_16793__1337 vssd1 vssd1 vccd1 vccd1 _16793__1337/HI net1337 sky130_fd_sc_hd__conb_1
XFILLER_0_206_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14959_ net1219 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XANTENNA__13473__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10287__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ net1064 _04170_ net1047 net959 vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12809__B _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16629_ clknet_leaf_94_wb_clk_i _02748_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13225__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09444__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] net765 net842 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\]
+ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16731__1359 vssd1 vssd1 vccd1 vccd1 net1359 _16731__1359/LO sky130_fd_sc_hd__conb_1
XFILLER_0_150_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13420__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09032_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\] net830 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a22o_1
XANTENNA__13199__Y _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold300 team_02_WB.instance_to_wrap.top.a1.row2\[41\] vssd1 vssd1 vccd1 vccd1 net1662
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 team_02_WB.instance_to_wrap.top.a1.row2\[10\] vssd1 vssd1 vccd1 vccd1 net1673
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12036__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold322 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] vssd1
+ vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold333 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold344 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 team_02_WB.instance_to_wrap.ramaddr\[31\] vssd1 vssd1 vccd1 vccd1 net1717
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold366 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold388 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout802 _04535_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_8
X_09934_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net804 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\]
+ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a221o_1
Xhold399 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1112_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 _04521_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
Xfanout824 _04512_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
Xfanout835 _04506_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__buf_4
XANTENNA__09904__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 _04359_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_2
XANTENNA__13375__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] net729 net713 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a22o_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 _04550_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_8
Xhold1000 team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1 vccd1 vccd1 net2362
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
XANTENNA_fanout572_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 _04538_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
Xhold1022 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net1484 net1041 net991 team_02_WB.instance_to_wrap.ramaddr\[15\] vssd1 vssd1
+ vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
X_09796_ _05306_ _05308_ _05310_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nor4_2
Xhold1044 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 team_02_WB.instance_to_wrap.top.a1.row2\[25\] vssd1 vssd1 vccd1 vccd1 net2417
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1066 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net846 _04363_ _04368_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__and3_4
Xhold1077 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 team_02_WB.instance_to_wrap.top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 net2461
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13391__A net2158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ _04305_ _04285_ _04290_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_64_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09683__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07629_ _03349_ _03350_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__nand2_1
XANTENNA__13216__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10640_ _04277_ net1059 net1060 vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__mux2_1
XANTENNA__08657__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09435__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ net424 net409 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12735__A _06943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ net240 net2445 net566 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ net1615 net984 net966 _02994_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ net1699 net353 net612 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XANTENNA__14950__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__A1 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net361 net1565 net464 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11785__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net398 _06630_ _06628_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_166_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15607__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07564__A team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15931_ clknet_leaf_29_wb_clk_i _02071_ _00739_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11054_ net1728 net265 net640 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
X_10005_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] net743 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15862_ clknet_leaf_21_wb_clk_i _02002_ _00670_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_199_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ net1205 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
XANTENNA_input19_X net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ clknet_leaf_0_wb_clk_i _01933_ _00601_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15757__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__A0 _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14744_ net1197 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
X_11956_ net294 net2225 net586 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XANTENNA__09674__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10907_ _06271_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__or2_1
X_14675_ net1073 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
X_11887_ net287 net2489 net486 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11025__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16414_ clknet_leaf_85_wb_clk_i _02549_ _01222_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _06348_ _06352_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
X_13626_ net1050 net1051 team_02_WB.instance_to_wrap.top.a1.row2\[12\] _03103_ vssd1
+ vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09426__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ clknet_leaf_124_wb_clk_i _02485_ _01153_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11233__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _05877_ net385 vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nor2_1
X_13557_ _03289_ net1049 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12508_ net240 net1898 net448 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__mux2_1
X_13488_ team_02_WB.START_ADDR_VAL_REG\[28\] net1070 net1004 vssd1 vssd1 vccd1 vccd1
+ net212 sky130_fd_sc_hd__a21o_1
X_16276_ clknet_leaf_14_wb_clk_i _02416_ _01084_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12439_ net352 net1964 net454 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
X_15227_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[18\]
+ _00040_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_117_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ net1157 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ net1204 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
X_15089_ net1072 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
X_07980_ _03670_ _03700_ _03702_ _03698_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_130_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16532__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ net525 _05165_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nor2_1
X_08601_ net96 net1579 net957 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
X_09581_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\] net733 net712 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__a22o_1
X_08532_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\] _04177_ vssd1 vssd1 vccd1
+ vccd1 _04218_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09665__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload92_A clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08463_ _04154_ _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09688__X _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ _04090_ _04093_ _04099_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_174_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout320_A _06936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10983__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09015_ net1058 _04297_ _04313_ net952 vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__and4b_4
XFILLER_0_103_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08928__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 _02584_ vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold141 net139 vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 team_02_WB.instance_to_wrap.ramstore\[27\] vssd1 vssd1 vccd1 vccd1 net1514
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13386__A team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold174 team_02_WB.START_ADDR_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_02_WB.instance_to_wrap.top.a1.row1\[123\] vssd1 vssd1 vccd1 vccd1 net1547
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 net116 vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _05422_ _05426_ _05430_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__or4_1
Xfanout643 _04452_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_4
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XANTENNA__16697__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_2
Xfanout676 _04412_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_4
X_09848_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] net806 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\]
+ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a221o_1
Xfanout687 _04399_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_8
Xfanout698 _04391_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\] net719 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_161_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11810_ net248 net2061 net590 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
X_12790_ _06698_ _06671_ _06670_ _06669_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__and4b_1
XFILLER_0_96_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09656__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11741_ net238 net2426 net596 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08864__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11672_ _04695_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nand2_1
X_14460_ net1192 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XANTENNA__08943__A _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13411_ _03018_ _03020_ _03021_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__or4_4
XFILLER_0_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__inv_2
X_14391_ net1207 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792__1336 vssd1 vssd1 vccd1 vccd1 _16792__1336/HI net1336 sky130_fd_sc_hd__conb_1
XFILLER_0_36_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16130_ clknet_leaf_120_wb_clk_i _02270_ _00938_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13342_ net2352 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[4\]
+ sky130_fd_sc_hd__and2_1
X_10554_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__inv_2
XANTENNA_input83_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__B2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16061_ clknet_leaf_11_wb_clk_i _02201_ _00869_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13273_ team_02_WB.instance_to_wrap.top.pc\[23\] net1053 _06618_ net935 vssd1 vssd1
+ vccd1 vccd1 _02986_ sky130_fd_sc_hd__a22o_1
X_10485_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09774__A _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ net1676 net284 net612 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
X_15012_ net1162 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10726__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ net278 net2462 net462 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
XANTENNA__12404__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _05983_ net664 _06117_ _06613_ _06614_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__o221a_1
X_12086_ net1689 net283 net583 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XANTENNA__11528__B _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09344__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ net424 _06547_ _06357_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a21oi_1
X_15914_ clknet_leaf_32_wb_clk_i _02054_ _00722_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_16730__1358 vssd1 vssd1 vccd1 vccd1 net1358 _16730__1358/LO sky130_fd_sc_hd__conb_1
X_15845_ clknet_leaf_28_wb_clk_i _01985_ _00653_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15016__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11439__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15776_ clknet_leaf_109_wb_clk_i _01916_ _00584_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12988_ team_02_WB.instance_to_wrap.top.pc\[9\] _05537_ _07507_ vssd1 vssd1 vccd1
+ vccd1 _07508_ sky130_fd_sc_hd__a21boi_1
X_14727_ net1174 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ net348 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\] net482 vssd1
+ vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XANTENNA__08855__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09949__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14658_ net1129 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16085__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ _03112_ _03127_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nor2_1
XANTENNA__11206__A2 _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14589_ net1207 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16328_ clknet_leaf_24_wb_clk_i _02468_ _01136_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09280__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16259_ clknet_leaf_10_wb_clk_i _02399_ _01067_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_11_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput213 net213 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_0_112_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09032__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12314__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07637__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _03651_ _03685_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10455__A_N _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] net756 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\]
+ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a221o_1
XANTENNA__13131__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07894_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__inv_2
XANTENNA__09886__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\] net826 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a22o_1
XANTENNA__16667__D _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__A1 _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _05061_ _05080_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nand2_1
XANTENNA__09099__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09638__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08515_ team_02_WB.instance_to_wrap.top.a1.data\[5\] net959 vssd1 vssd1 vccd1 vccd1
+ _04205_ sky130_fd_sc_hd__or2_1
XFILLER_0_195_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09495_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] net702 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a22o_1
XANTENNA__08846__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16428__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08446_ _04130_ _04139_ _04142_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_176_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08377_ _04081_ _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_A _04389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12158__A0 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10270_ _04326_ _04492_ _05786_ net650 vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12224__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10184__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__B2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _07226_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_6
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _07222_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_21_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout473 _07208_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_8
X_13960_ net1167 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
Xfanout484 _07200_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09877__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout495 _06252_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_2
XFILLER_0_198_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11635__Y _07122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ _07361_ _07430_ _07362_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o21a_1
X_13891_ net1246 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
X_15630_ clknet_leaf_61_wb_clk_i _01770_ _00438_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _04494_ _04886_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09629__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15561_ clknet_leaf_111_wb_clk_i _01701_ _00369_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12773_ net546 _06118_ _06402_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__and4_1
XFILLER_0_185_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08837__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14512_ net1236 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11724_ net315 net2065 net602 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15492_ clknet_leaf_36_wb_clk_i _01632_ _00300_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11655_ _05649_ _05922_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_30_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14443_ net1098 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12397__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10606_ _04461_ _06114_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14374_ net1204 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
X_11586_ _05910_ _06000_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09801__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16113_ clknet_leaf_0_wb_clk_i _02253_ _00921_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10537_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__inv_2
X_13325_ net1620 _03010_ _03012_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12149__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap618 _07215_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ clknet_leaf_2_wb_clk_i _02184_ _00852_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10468_ _05212_ _05977_ _05980_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__or4_1
X_13256_ team_02_WB.instance_to_wrap.top.pc\[29\] net1055 net934 _02974_ vssd1 vssd1
+ vccd1 vccd1 _02975_ sky130_fd_sc_hd__a22o_1
XANTENNA__08612__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12207_ net363 net2452 net576 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
XANTENNA__12134__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _07495_ _07498_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__xor2_1
X_10399_ _05691_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nor2_2
X_12138_ net358 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\] net467 vssd1
+ vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11973__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ net339 net2443 net473 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09868__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15828_ clknet_leaf_114_wb_clk_i _01968_ _00636_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15759_ clknet_leaf_48_wb_clk_i _01899_ _00567_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08300_ _03985_ _04010_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09280_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\] net730 net715 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08231_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _03840_ _03847_ net227 _03841_ _03802_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09253__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__X _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08093_ _03759_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11__f_wb_clk_i_X clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload50 clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_16
Xclkload61 clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__inv_16
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08522__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload72 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload72/X sky130_fd_sc_hd__clkbuf_8
Xclkload83 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload94 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload94/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12044__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ net944 _04503_ _04505_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout485_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _03666_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_145_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11115__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09859__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16791__1335 vssd1 vssd1 vccd1 vccd1 _16791__1335/HI net1335 sky130_fd_sc_hd__conb_1
XFILLER_0_208_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07877_ _03574_ _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout652_A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09616_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\] net766 _05130_ _05132_
+ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_178_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] net834 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\]
+ _05063_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a221o_1
XANTENNA__08819__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1182_X net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ _04970_ _04991_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08429_ _04128_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__or2_1
XANTENNA__12219__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15968__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11440_ net1882 net319 net637 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
Xclkload0 clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__inv_6
XFILLER_0_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11371_ _06772_ _06869_ net396 vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\] net922 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a22o_1
X_13110_ _07371_ _07419_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__nor2_1
X_14090_ net1118 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_189_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13041_ _07355_ _07437_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__xnor2_1
X_10253_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\] net746 _05767_ _05768_
+ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10157__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\] net802 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\]
+ _05700_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__a221o_1
Xfanout1202 net1265 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_2
XANTENNA_input46_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1213 net1218 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
Xfanout1224 net1227 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_4
XANTENNA__11793__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1246 net1248 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_208_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1257 net1262 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_4
X_14992_ net1155 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08668__A team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 _06657_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_1
XANTENNA__07572__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16731_ net1359 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xfanout292 _06791_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
X_13943_ net1249 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16662_ clknet_leaf_93_wb_clk_i _02781_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13874_ net1164 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15613_ clknet_leaf_13_wb_clk_i _01753_ _00421_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12825_ _03319_ _07340_ _07341_ _04172_ _03317_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__o32a_1
X_16593_ clknet_leaf_96_wb_clk_i _02712_ _01386_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15544_ clknet_leaf_122_wb_clk_i _01684_ _00352_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12756_ _05647_ _05691_ _07278_ _07279_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__or4_1
XANTENNA__08607__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_X clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_154_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ net237 net1985 net600 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XANTENNA__12129__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15475_ clknet_leaf_58_wb_clk_i _01615_ _00283_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12687_ net292 net1989 net431 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__mux2_1
X_14426_ net1097 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11638_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] _04347_ net953 _07124_ vssd1
+ vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11968__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ net1224 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11569_ net418 _06694_ _06898_ net376 _07055_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16123__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold718 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ net1640 net984 net966 _03003_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__a22o_1
Xhold729 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13468__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14288_ net1232 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
X_16027_ clknet_leaf_32_wb_clk_i _02167_ _00835_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13239_ _02953_ _02958_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__nand2_1
XANTENNA__09002__A3 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10148__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _03515_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08761__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08780_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] net769 net677 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\]
+ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10901__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire620_A _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07731_ _03386_ _03411_ _03418_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09026__X _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10620__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08297__B _03746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07662_ _03347_ _03379_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_0_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10320__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\] net751 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07593_ team_02_WB.instance_to_wrap.top.a1.state\[1\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__or3_1
XFILLER_0_177_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09332_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] net901 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__a22o_1
XANTENNA__09474__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_173_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12039__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08214_ _03901_ _03921_ _03927_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09226__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09194_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] net730 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11878__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _03829_ _03836_ net227 vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1142_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13378__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03787_ _03762_ vssd1 vssd1
+ vccd1 vccd1 _03797_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10139__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_X net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\] vssd1 vssd1 vccd1 vccd1
+ net1374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13394__A net2615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\] vssd1 vssd1 vccd1 vccd1
+ net1385 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 team_02_WB.instance_to_wrap.ramstore\[14\] vssd1 vssd1 vccd1 vccd1 net1396
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net1063 net1062 _04267_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a21oi_1
Xhold45 team_02_WB.instance_to_wrap.ramstore\[26\] vssd1 vssd1 vccd1 vccd1 net1407
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _02563_ vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_02_WB.instance_to_wrap.ramaddr\[3\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07929_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03648_ _03649_ _03650_ vssd1
+ vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__o211a_1
XANTENNA__11639__A2 _07122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold78 _02599_ vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15382__Q team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 team_02_WB.instance_to_wrap.ramstore\[4\] vssd1 vssd1 vccd1 vccd1 net1451
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ _06355_ _06452_ net656 vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_203_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ _06384_ _06385_ net394 vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15790__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12610_ net2390 net255 net553 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XANTENNA__11642__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input100_A wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ team_02_WB.instance_to_wrap.top.a1.row2\[41\] _03123_ _03125_ team_02_WB.instance_to_wrap.top.a1.row2\[33\]
+ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a221o_1
XANTENNA__09465__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ net242 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\] net444 vssd1
+ vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14953__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15260_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[19\]
+ _00073_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ net351 net2241 net450 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ net1132 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XANTENNA__11788__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ _06868_ _06919_ net370 vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15191_ net1145 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10378__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__B team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _06354_ _06853_ _06850_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__o21bai_2
XANTENNA__07567__A team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14142_ net1188 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10305_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] net713 _05820_ _05821_
+ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a211o_1
XANTENNA__13316__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14073_ net1089 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
X_11285_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] net494 _06787_ _04263_ net496
+ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10236_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] net802 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a221o_1
X_13024_ net1026 _07543_ net1024 team_02_WB.instance_to_wrap.top.pc\[31\] vssd1 vssd1
+ vccd1 vccd1 _01512_ sky130_fd_sc_hd__a2bb2o_1
Xfanout1010 _03314_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_2
XANTENNA__12412__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1032 net1033 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__buf_2
X_10167_ _05677_ _05679_ _05681_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or4_1
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_2
Xfanout1054 net1056 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13221__A1_N net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_4
XFILLER_0_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1087 net1094 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_4
X_14975_ net1160 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
X_10098_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\] net714 _05612_ _05613_
+ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__a2111o_1
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16714_ net1273 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13926_ net1234 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10302__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16645_ clknet_leaf_93_wb_clk_i _02764_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13857_ net1148 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12808_ _07330_ _07331_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__and2b_2
XANTENNA__09456__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16576_ clknet_leaf_93_wb_clk_i _00002_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13788_ net2419 _03276_ net961 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__o21ai_1
X_15527_ clknet_leaf_42_wb_clk_i _01667_ _00335_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12739_ net795 _06108_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ clknet_leaf_119_wb_clk_i _01598_ _00266_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16790__1334 vssd1 vssd1 vccd1 vccd1 _16790__1334/HI net1334 sky130_fd_sc_hd__conb_1
X_14409_ net1221 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ clknet_leaf_13_wb_clk_i _01529_ _00197_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10369__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold504 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10615__B _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold537 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__inv_2
Xhold559 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09692__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15663__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ net13 net1032 net988 net1601 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
X_09881_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\] net709 _05394_ _05395_
+ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_51_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12830__B _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] _03301_ team_02_WB.instance_to_wrap.wb.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__and3b_4
XANTENNA__12322__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10631__A team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1204 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1237 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\] net721 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__a22o_1
Xhold1259 team_02_WB.instance_to_wrap.top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 net2621
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07714_ _03431_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__and2_1
XANTENNA__13942__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08595__X _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ net1062 _04309_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12829__Y _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _03364_ _03365_ _03366_ vssd1
+ vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout350_A _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__and2b_1
XANTENNA__09447__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\] net783 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09246_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\] net828 net812 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\]
+ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_153_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09177_ _04656_ _04661_ _04671_ _04692_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_153_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13546__A2 _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ _03846_ _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15377__Q team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1253_X net2615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08059_ _03736_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_101_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11070_ net381 _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] net896 net943 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a22o_1
Xinput102 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12232__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ net1113 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XANTENNA__09686__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11972_ net353 net2450 net584 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09150__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03227_ _03229_ vssd1
+ vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__o21a_1
X_10923_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14691_ net1136 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16430_ clknet_leaf_61_wb_clk_i net1460 _01238_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ team_02_WB.instance_to_wrap.top.a1.row1\[15\] _03113_ _03109_ vssd1 vssd1
+ vccd1 vccd1 _03190_ sky130_fd_sc_hd__o21a_1
XANTENNA__09113__Y _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10854_ _06131_ net653 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] net496
+ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_4_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ clknet_leaf_113_wb_clk_i _02501_ _01169_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13573_ _03107_ _03127_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nor2_1
XANTENNA__15536__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10785_ _05440_ net404 vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15312_ clknet_leaf_44_wb_clk_i _01455_ _00125_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12524_ net308 net2330 net447 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16292_ clknet_leaf_36_wb_clk_i _02432_ _01100_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15243_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[2\]
+ _00056_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12455_ net285 net2562 net450 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__mux2_1
XANTENNA__12407__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ _05378_ net660 net659 _05379_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a22o_1
X_15174_ net1142 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12386_ net278 net2262 net458 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14125_ net1126 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XANTENNA__08964__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11337_ _06836_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__or2_1
XANTENNA__08620__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ net1111 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
X_11268_ _05103_ net386 _06089_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__o21ai_1
X_13007_ _07458_ _07526_ _07459_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__o21bai_1
X_10219_ net422 net502 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__nor2_1
XANTENNA__12142__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10451__A _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ _04469_ _06687_ _06704_ net671 _06703_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__a221o_4
XANTENNA__14858__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11981__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14958_ net1076 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XANTENNA__09677__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16311__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09141__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13175__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ net1261 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14889_ net1217 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
X_16628_ clknet_leaf_94_wb_clk_i _02747_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13225__B2 _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10039__A1 _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16559_ clknet_leaf_87_wb_clk_i _02683_ _01366_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08101__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\] net681 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] net818 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12317__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09974__X _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13113__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold323 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_02_WB.instance_to_wrap.ramload\[24\] vssd1 vssd1 vccd1 vccd1 net1696
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold345 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold378 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\] net902 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a22o_1
Xhold389 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 _04535_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08530__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout814 _04521_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_209_Left_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout825 _04512_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12052__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__inv_2
Xfanout847 _04358_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_2
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_181_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1105_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 _04541_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_4
Xhold1012 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ net113 net1045 net992 net1482 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1023 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\] net740 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a221o_1
Xhold1034 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout565_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1045 team_02_WB.instance_to_wrap.top.pad.keyCode\[2\] vssd1 vssd1 vccd1 vccd1
+ net2407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11891__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_02_WB.instance_to_wrap.top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 net2429
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _04302_ net846 _04365_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__and3_1
XANTENNA__09668__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1078 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 team_02_WB.instance_to_wrap.top.a1.row1\[121\] vssd1 vssd1 vccd1 vccd1 net2451
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout732_A _04381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07628_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] _03348_ vssd1 vssd1 vccd1
+ vccd1 _03351_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13216__B2 _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[3\] vssd1 vssd1 vccd1 vccd1
+ _03300_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1262_X net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10570_ net419 net413 vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\] net842 _04740_ _04742_
+ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12227__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ net1806 net364 net612 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XANTENNA__09199__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_86_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13847__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ net342 net1761 net463 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
XANTENNA__08946__A2 _04339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11122_ _06576_ _06629_ net371 vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__mux2_1
Xhold890 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13152__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11053_ net947 _06556_ _06563_ net606 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__o211a_2
X_15930_ clknet_leaf_50_wb_clk_i _02070_ _00738_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10271__A _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\] net788 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09371__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ clknet_leaf_31_wb_clk_i _02001_ _00669_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_199_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ net1193 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_199_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09659__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15792_ clknet_leaf_30_wb_clk_i _01932_ _00600_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10269__A1 _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ net1207 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11955_ net286 net1970 net584 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10906_ team_02_WB.instance_to_wrap.top.pc\[29\] _06270_ vssd1 vssd1 vccd1 vccd1
+ _06421_ sky130_fd_sc_hd__nor2_1
X_14674_ net1178 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
X_11886_ net274 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\] net488 vssd1
+ vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__mux2_1
XANTENNA__08882__B2 net2158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16413_ clknet_leaf_99_wb_clk_i _02548_ _01221_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ net1405 net962 _03176_ net1067 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16344_ clknet_leaf_114_wb_clk_i _02484_ _01152_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ net1051 _03290_ _03109_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10768_ _04611_ _06033_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ net641 _07203_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__nand2_4
XFILLER_0_81_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12137__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16275_ clknet_leaf_57_wb_clk_i _02415_ _01083_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13487_ team_02_WB.START_ADDR_VAL_REG\[27\] net1071 net1005 vssd1 vssd1 vccd1 vccd1
+ net211 sky130_fd_sc_hd__a21o_1
X_10699_ team_02_WB.instance_to_wrap.top.pc\[17\] _06190_ vssd1 vssd1 vccd1 vccd1
+ _06216_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15226_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[17\]
+ _00039_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12438_ net364 net1743 net454 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11976__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10880__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15157_ net1159 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
X_12369_ net343 net2076 net561 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14108_ net1201 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
X_15088_ net1078 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ net1207 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XANTENNA__09018__Y _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ _04249_ _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nand2_4
XFILLER_0_207_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09580_ _05085_ _05089_ _05093_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or4_1
XANTENNA__12600__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ team_02_WB.instance_to_wrap.top.a1.data\[1\] net959 vssd1 vssd1 vccd1 vccd1
+ _04217_ sky130_fd_sc_hd__or2_1
XANTENNA__11457__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08462_ _04158_ _04160_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1
+ vccd1 vccd1 _04164_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_46_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08393_ _04082_ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12836__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09822__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12047__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1055_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09014_ _04297_ _04313_ net945 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11886__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold120 team_02_WB.instance_to_wrap.ramaddr\[16\] vssd1 vssd1 vccd1 vccd1 net1482
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold131 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold142 _02562_ vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _02589_ vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13386__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 team_02_WB.instance_to_wrap.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 net1537
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 team_02_WB.START_ADDR_VAL_REG\[1\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout600 _07189_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_57_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold197 _02613_ vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] net777 _05431_ _05432_
+ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a211o_1
XANTENNA_hold1049_X net2411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net656 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_148_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09353__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_2
Xfanout677 net680 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_8
X_09847_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] net908 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a22o_1
Xfanout688 _04399_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XANTENNA__14498__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12510__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_161_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09105__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11448__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] net931 vssd1 vssd1 vccd1
+ vccd1 _04358_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11740_ net245 net2623 net598 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
XANTENNA__10120__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ _04569_ _04611_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08943__B _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13410_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__or4b_1
X_10622_ net551 _06128_ _06138_ _06126_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14390_ net1106 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09813__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13341_ team_02_WB.instance_to_wrap.ramload\[3\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[3\] sky130_fd_sc_hd__and2_1
X_10553_ _06054_ _06069_ net412 vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10266__A _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10974__A2 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16060_ clknet_leaf_16_wb_clk_i _02200_ _00868_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input76_A wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ net1612 net982 net964 _02985_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _05907_ _06000_ _05908_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11796__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ net1160 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
X_12223_ net2530 net272 net615 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XANTENNA__10187__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ net280 net2177 net464 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
XANTENNA__09592__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__X _03746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _04907_ _06113_ _06116_ _04908_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o22a_1
X_12085_ net2474 net270 net583 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
X_11036_ net409 _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__nor2_1
X_15913_ clknet_leaf_115_wb_clk_i _02053_ _00721_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11384__X _06883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15844_ clknet_leaf_35_wb_clk_i _01984_ _00652_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12420__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14201__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15775_ clknet_leaf_59_wb_clk_i _01915_ _00583_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12987_ _07505_ _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14726_ net1218 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11938_ net350 net2420 net482 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XANTENNA__10111__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ net1262 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
XANTENNA__09949__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ net364 net1907 net490 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13608_ _03115_ _03120_ _03116_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a21o_1
XANTENNA__09804__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14588_ net1192 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16327_ clknet_leaf_38_wb_clk_i _02467_ _01135_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13539_ team_02_WB.instance_to_wrap.top.edg2.button_i _03074_ _03083_ _03087_ vssd1
+ vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_41_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15254__CLK clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16258_ clknet_leaf_117_wb_clk_i _02398_ _01066_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15209_ clknet_leaf_97_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[0\]
+ _00022_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] sky130_fd_sc_hd__dfrtp_4
Xoutput203 net203 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput214 net214 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
X_16189_ clknet_leaf_12_wb_clk_i _02329_ _00997_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10178__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10904__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09583__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__Y _05488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03648_ _03670_ _03672_ vssd1
+ vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__a2bb2o_1
X_09701_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\] net774 net770 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a22o_1
XANTENNA__09335__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ _03580_ _03606_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__xnor2_1
X_09632_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] net805 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ _05148_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a221o_1
XANTENNA__12330__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09563_ net970 net630 net544 vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout263_A _06595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16739__1284 vssd1 vssd1 vccd1 vccd1 _16739__1284/HI net1284 sky130_fd_sc_hd__conb_1
XFILLER_0_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ _04204_ net1621 _04186_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
XANTENNA__13950__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] net749 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\]
+ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a221o_1
XANTENNA__10102__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10653__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ _04141_ _04146_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout430_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1172_A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ net1748 net1006 net981 _04086_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08074__A2 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_A _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12505__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09574__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _07229_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_8
Xfanout441 _07226_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09326__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_6
Xfanout463 _07213_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 _07206_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_6
Xfanout485 _07200_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_4
X_12910_ _04928_ _06177_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__a21o_1
Xfanout496 net497 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
XANTENNA__12240__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15117__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ net1253 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10341__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12841_ _04494_ _04886_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_17_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15560_ clknet_leaf_11_wb_clk_i _01700_ _00368_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12772_ _06579_ _06606_ net381 vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_169_Left_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14511_ net1219 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_11723_ net306 net2374 net603 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15491_ clknet_leaf_27_wb_clk_i _01631_ _00299_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15277__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14442_ net1117 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
X_11654_ _05468_ _07139_ _06011_ _06956_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_71_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _04461_ _06114_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__nor2_4
XFILLER_0_154_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14373_ net1117 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
X_11585_ net418 _06726_ _06921_ net376 _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__a221o_2
X_16112_ clknet_leaf_23_wb_clk_i _02252_ _00920_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13324_ _04169_ _03010_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10536_ _06044_ _06052_ net395 vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16043_ clknet_leaf_15_wb_clk_i _02183_ _00851_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13255_ _02965_ _02973_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ _04951_ _05983_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_178_Left_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12415__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12206_ net354 net2020 net578 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13186_ _07389_ _07393_ _07394_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_57_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10398_ net504 _05690_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__and2_1
X_12137_ net342 net2351 net468 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09317__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12068_ net333 net2314 net470 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12150__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ net1858 net258 net637 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XANTENNA__10332__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15827_ clknet_leaf_59_wb_clk_i _01967_ _00635_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15758_ clknet_leaf_47_wb_clk_i _01898_ _00566_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14709_ net1242 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
X_15689_ clknet_leaf_110_wb_clk_i _01829_ _00497_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08230_ _03935_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10618__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08161_ _03840_ _03847_ net227 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08092_ _03771_ _03776_ _03781_ _03787_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12833__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload40 clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__clkinv_2
Xclkload51 clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_12
XANTENNA__12325__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload62 clknet_leaf_86_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_12
Xclkload73 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload73/X sky130_fd_sc_hd__clkbuf_8
Xclkload84 clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload84/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09556__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload95 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_6
XANTENNA__08104__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13945__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11362__A1_N net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ net945 _04507_ _04509_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__and3_4
XANTENNA__09308__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _03626_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_145_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ _03596_ _03597_ _03586_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10323__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11520__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\] net718 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\]
+ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09546_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\] net871 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a22o_1
XANTENNA__08774__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _04970_ _04992_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout812_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__A _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1175_X net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08428_ net1652 net1006 net981 _04134_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ net2282 net1006 net980 _04070_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_210_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09795__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ _06818_ _06868_ net370 vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11199__X _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10321_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] net828 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\]
+ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__a221o_1
XANTENNA__12235__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__A _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11339__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09547__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ _07535_ _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__xnor2_1
X_10252_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] net775 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a22o_1
X_10183_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] net921 net885 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__a22o_1
Xfanout1203 net1206 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 net1218 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
X_16759__1303 vssd1 vssd1 vccd1 vccd1 _16759__1303/HI net1303 sky130_fd_sc_hd__conb_1
XFILLER_0_206_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1225 net1227 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_2
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14991_ net1135 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1247 net1248 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1258 net1259 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
Xfanout260 _06530_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16075__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11106__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 _06626_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
XANTENNA__08668__B team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_2
X_16730_ net1358 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
X_13942_ net1249 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
Xfanout293 _06791_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_199_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09180__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ clknet_leaf_93_wb_clk_i _02780_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13873_ net1165 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ clknet_leaf_17_wb_clk_i _01752_ _00420_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12824_ team_02_WB.instance_to_wrap.top.a1.state\[1\] _07343_ _07345_ _07341_ vssd1
+ vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__o22a_1
X_16592_ clknet_leaf_90_wb_clk_i _02711_ _01385_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08684__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15543_ clknet_leaf_122_wb_clk_i _01683_ _00351_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ _05736_ _05783_ _05829_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_201_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11314__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ net244 net2441 net602 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XANTENNA__10093__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15474_ clknet_leaf_54_wb_clk_i _01614_ _00282_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12686_ net286 net1875 net430 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__mux2_1
XANTENNA__08971__X _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14425_ net1097 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ net1001 net995 _07123_ team_02_WB.instance_to_wrap.top.pc\[1\] vssd1 vssd1
+ vccd1 vccd1 _07124_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11042__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11042__B2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09786__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ net1239 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
X_11568_ _05738_ _06001_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__xor2_1
XANTENNA__08623__S _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold708 net107 vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ team_02_WB.instance_to_wrap.top.pc\[6\] net1054 _07026_ net933 vssd1 vssd1
+ vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_1
X_10519_ net669 _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__nor2_1
Xhold719 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_1
XANTENNA__10454__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14287_ net1220 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
XANTENNA__12145__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11499_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _06833_ _06837_ _06992_ vssd1
+ vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16026_ clknet_leaf_19_wb_clk_i _02166_ _00834_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09538__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ team_02_WB.instance_to_wrap.top.ru.next_write_i _00006_ vssd1 vssd1 vccd1
+ vccd1 _02959_ sky130_fd_sc_hd__nor2_4
X_16738__1283 vssd1 vssd1 vccd1 vccd1 _16738__1283/HI net1283 sky130_fd_sc_hd__conb_1
XANTENNA__11984__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16418__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13169_ net1026 _02931_ net1023 team_02_WB.instance_to_wrap.top.pc\[7\] vssd1 vssd1
+ vccd1 vccd1 _01488_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13484__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10901__B _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _03443_ _03447_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09171__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07661_ _03344_ _03370_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09710__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] net776 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\]
+ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07592_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] _03316_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 _03317_
+ sky130_fd_sc_hd__or4b_4
X_09331_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\] net835 net831 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09474__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _04777_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08213_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09193_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\] net715 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a22o_1
XANTENNA__12844__A _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08144_ _03829_ _03835_ net227 vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11584__A2 _06998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03787_ vssd1 vssd1 vccd1
+ vccd1 _03796_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12055__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1135_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09529__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16098__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A _07192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 team_02_WB.instance_to_wrap.ramaddr\[30\] vssd1 vssd1 vccd1 vccd1 net1375
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_02_WB.instance_to_wrap.ramstore\[30\] vssd1 vssd1 vccd1 vccd1 net1386
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _04491_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and2_2
Xhold35 _02576_ vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 _02588_ vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12297__A0 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07928_ _03649_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nand2_1
Xhold57 team_02_WB.instance_to_wrap.top.a1.data\[4\] vssd1 vssd1 vccd1 vccd1 net1419
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _02597_ vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_02_WB.instance_to_wrap.ramstore\[24\] vssd1 vssd1 vccd1 vccd1 net1441
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10847__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__B2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _03540_ _03544_ _03545_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ _06058_ _06063_ net369 vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09529_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] net731 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ net641 _07205_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__nand2_8
XANTENNA__10075__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ net362 net2624 net450 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__mux2_1
XANTENNA__08951__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210_ net1129 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_193_Right_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11422_ net517 _05901_ _06061_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15190_ net1141 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XANTENNA__09768__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__A1 _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08670__C team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ net1203 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ _06358_ _06638_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_111_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10304_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\] net753 net729 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14072_ net1196 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11284_ _06786_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__inv_2
X_13023_ _06273_ net233 _07443_ net977 _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__o221a_1
X_10235_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] net834 net814 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1000 _04264_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
Xfanout1022 _00012_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09940__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1033 _04429_ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_2
X_10166_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\] net829 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a221o_1
Xfanout1044 net1046 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1068 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
Xfanout1077 net1101 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_4
Xfanout1088 net1094 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_2
X_10097_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\] net734 net720 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a22o_1
X_14974_ net1164 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_4
X_16713_ net1272 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13925_ net1244 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload4_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__X _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16644_ clknet_leaf_92_wb_clk_i _02763_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13856_ net1147 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08618__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _07234_ _07231_ _06124_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10449__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13787_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ _03275_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__and3_1
X_16575_ clknet_leaf_92_wb_clk_i _00001_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10999_ _06447_ _06510_ net372 vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__mux2_1
XANTENNA__13252__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ net380 _06579_ _06518_ _06484_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15526_ clknet_leaf_6_wb_clk_i _01666_ _00334_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11979__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15457_ clknet_leaf_101_wb_clk_i _01597_ _00265_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12669_ net364 net2091 net434 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14408_ net1115 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XANTENNA__09759__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15388_ clknet_leaf_19_wb_clk_i _01528_ _00196_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08967__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14339_ net1132 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold505 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap224 _03949_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_1
Xhold516 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold549 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08719__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16009_ clknet_leaf_116_wb_clk_i _02149_ _00817_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_08900_ net24 net1033 net988 team_02_WB.instance_to_wrap.ramload\[2\] vssd1 vssd1
+ vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
X_09880_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\] net705 _05396_ vssd1
+ vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a21o_1
XANTENNA__12603__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ net1569 net1038 net990 team_02_WB.instance_to_wrap.ramaddr\[0\] vssd1 vssd1
+ vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XANTENNA__09931__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1205 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10631__B _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1216 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15958__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1227 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ _04296_ net846 _04363_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__and3_2
Xhold1238 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10829__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03432_ _03433_ _03434_ vssd1
+ vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a2bb2o_1
X_08693_ _04294_ _04319_ _04321_ _04310_ _04317_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o311a_1
XANTENNA__13491__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07644_ _03365_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ net2579 net189 _00017_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout343_A _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1085_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\] net747 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a22o_1
XANTENNA__11254__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10057__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09998__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11889__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\] net878 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16758__1302 vssd1 vssd1 vccd1 vccd1 _16758__1302/HI net1302 sky130_fd_sc_hd__conb_1
XFILLER_0_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1252_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09176_ net542 _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08958__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ _03803_ _03841_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1040_X net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1138_X net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15488__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08058_ _03757_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__A _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10020_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_168_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09922__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput103 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09135__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11971_ net365 net1947 net584 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
X_13710_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03227_ net1139 vssd1
+ vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a21oi_1
X_10922_ net408 _06435_ _06434_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10296__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14690_ net1130 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13641_ _03167_ _03181_ _03188_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__or3_1
X_10853_ net999 _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_197_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10048__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16360_ clknet_leaf_16_wb_clk_i _02500_ _01168_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13572_ _03104_ _03115_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nand2_1
XANTENNA__09989__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ _05489_ net385 vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15311_ clknet_leaf_61_wb_clk_i _01454_ _00124_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11799__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ net302 net2254 net448 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__mux2_1
X_16291_ clknet_leaf_26_wb_clk_i _02431_ _01099_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15242_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[1\]
+ _00055_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12454_ net273 net2384 net452 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08949__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ net416 _06438_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15173_ net1143 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
X_12385_ net282 net2024 net460 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14124_ net1209 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11336_ net848 net953 net497 vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__o21a_2
XANTENNA__12931__B _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14055_ net1180 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
X_11267_ net374 _06535_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12423__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09374__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ team_02_WB.instance_to_wrap.top.pc\[21\] _06184_ _07525_ vssd1 vssd1 vccd1
+ vccd1 _07526_ sky130_fd_sc_hd__a21oi_1
X_10218_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] net780 _05728_ _05733_
+ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a2111oi_1
XPHY_EDGE_ROW_105_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10845__A2_N net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09913__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ _05041_ _06600_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__xnor2_1
X_10149_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] net738 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09126__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14957_ net1121 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XANTENNA__13473__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10287__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ net1248 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XANTENNA__09304__Y _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14888_ net1105 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16627_ clknet_leaf_94_wb_clk_i _02746_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ net1155 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_114_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16558_ clknet_leaf_87_wb_clk_i _02682_ _01365_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[109\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ clknet_leaf_31_wb_clk_i _01649_ _00317_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16489_ clknet_leaf_66_wb_clk_i net1376 _01297_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09030_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] net928 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold302 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12841__B _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold368 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\] net882 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12333__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold379 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_123_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 _04534_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09365__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout815 _04521_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_4
Xfanout826 _04512_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_8
X_09863_ _05378_ _05379_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nand2b_1
Xfanout837 _04470_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
XANTENNA__09904__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 _04325_ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_2
XANTENNA__10361__B _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _04544_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_181_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ net1516 net1040 net991 team_02_WB.instance_to_wrap.ramaddr\[17\] vssd1 vssd1
+ vccd1 vccd1 _02611_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_181_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\] net736 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a22o_1
Xhold1024 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1035 team_02_WB.instance_to_wrap.ramload\[0\] vssd1 vssd1 vccd1 vccd1 net2397
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09117__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1057 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\] vssd1
+ vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _04358_ _04365_ _04370_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__and3_1
Xhold1068 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10278__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _04262_ _04293_ _04294_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_200_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07627_ _03324_ _03327_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1
+ vccd1 vccd1 _03350_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_132_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13216__A2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07558_ team_02_WB.instance_to_wrap.top.edg2.flip2 vssd1 vssd1 vccd1 vccd1 _03299_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_119_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10817__A _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1255_X net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] net777 _04743_ _04744_
+ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13220__A1_N _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09159_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\] net891 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\]
+ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10202__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ net340 net1914 net463 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_141_Left_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _06320_ _06339_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold880 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _06557_ _06562_ _06561_ _06558_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a211o_1
X_10003_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] net776 _05517_ _05519_
+ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a211o_1
X_15860_ clknet_leaf_14_wb_clk_i _02000_ _00668_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09108__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14811_ net1077 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15791_ clknet_leaf_41_wb_clk_i _01931_ _00599_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ net275 net1798 net586 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_150_Left_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14742_ net1107 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _06134_ net652 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] net496
+ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a221o_1
X_14673_ net1226 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net289 net2302 net489 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13624_ team_02_WB.instance_to_wrap.top.a1.row2\[27\] _03118_ _03169_ _03170_ _03175_
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__a2111o_1
X_16412_ clknet_leaf_80_wb_clk_i _02547_ _01220_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10836_ _06349_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16343_ clknet_leaf_122_wb_clk_i _02483_ _01151_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13555_ net1051 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03109_ vssd1
+ vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__and3_1
X_10767_ _04611_ _05959_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__xor2_1
XANTENNA__12418__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ net346 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\] net556 vssd1
+ vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__mux2_1
X_16274_ clknet_leaf_54_wb_clk_i _02414_ _01082_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13486_ team_02_WB.START_ADDR_VAL_REG\[26\] net1071 net1005 vssd1 vssd1 vccd1 vccd1
+ net210 sky130_fd_sc_hd__a21o_1
XFILLER_0_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ team_02_WB.instance_to_wrap.top.pc\[16\] _06192_ _06214_ vssd1 vssd1 vccd1
+ vccd1 _06215_ sky130_fd_sc_hd__a21o_1
XANTENNA__10446__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15225_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[16\]
+ _00038_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_12437_ net356 net2392 net456 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09595__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15156_ net1159 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
X_12368_ net339 net2157 net560 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14107_ net1085 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11319_ _06715_ _06819_ net400 vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12153__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15087_ net1079 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
X_12299_ net326 net2394 net569 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14038_ net1083 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XFILLER_0_180_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11992__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16757__1301 vssd1 vssd1 vccd1 vccd1 _16757__1301/HI net1301 sky130_fd_sc_hd__conb_1
X_15989_ clknet_leaf_40_wb_clk_i _02129_ _00797_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11293__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _04216_ net1581 net849 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
XANTENNA__11457__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08461_ net1602 net1008 net981 _04163_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08392_ _04090_ _04092_ _04099_ _04088_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__o31a_1
XANTENNA__10680__A2 _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12836__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12328__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ net1058 _04528_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__nor2_8
XANTENNA__13948__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold110 team_02_WB.instance_to_wrap.ramaddr\[27\] vssd1 vssd1 vccd1 vccd1 net1472
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _02610_ vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold132 team_02_WB.instance_to_wrap.top.a1.row1\[104\] vssd1 vssd1 vccd1 vccd1 net1494
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 team_02_WB.instance_to_wrap.top.pad.button_control.noisy vssd1 vssd1 vccd1
+ vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold154 net114 vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net1527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12063__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold176 _02571_ vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 _07189_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_4
Xhold187 net122 vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 team_02_WB.instance_to_wrap.top.a1.row2\[2\] vssd1 vssd1 vccd1 vccd1 net1560
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _07215_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_6
X_09915_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\] net709 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout656 _06123_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
Xfanout667 _06038_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_4
X_09846_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\] net811 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\]
+ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a221o_1
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_8
Xfanout689 _04397_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _05292_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08728_ team_02_WB.instance_to_wrap.top.i_ready net1001 net790 net551 vssd1 vssd1
+ vccd1 vccd1 _04357_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ net1061 net1059 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11670_ _05987_ _07155_ _07150_ _05986_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10621_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net995 vssd1 vssd1 vccd1
+ vccd1 _06138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10547__A _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13340_ team_02_WB.instance_to_wrap.ramload\[2\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[2\] sky130_fd_sc_hd__and2_1
X_10552_ _06060_ _06068_ net393 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__mux2_1
XANTENNA__11081__C1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13271_ team_02_WB.instance_to_wrap.top.pc\[24\] net1055 _06588_ net933 vssd1 vssd1
+ vccd1 vccd1 _02985_ sky130_fd_sc_hd__a22o_1
X_10483_ net408 net498 _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__o21ai_1
X_15010_ net1135 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
XANTENNA__09577__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ net1713 net288 net613 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
XANTENNA__16301__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input69_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ net271 net1768 net465 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ net380 _06606_ _06357_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09329__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__B2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ net2612 net264 net583 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XANTENNA__11136__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14689__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _05809_ _06350_ _06400_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__a31o_1
X_15912_ clknet_leaf_24_wb_clk_i _02052_ _00720_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11687__A1 _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15843_ clknet_leaf_27_wb_clk_i _01983_ _00651_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11439__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15774_ clknet_leaf_5_wb_clk_i _01914_ _00582_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12986_ team_02_WB.instance_to_wrap.top.pc\[9\] _05536_ vssd1 vssd1 vccd1 vccd1 _07506_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09501__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14725_ net1176 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
X_11937_ net362 net2463 net482 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XANTENNA__08855__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11868_ net357 net2172 net492 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
XANTENNA__08626__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14656_ net1103 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ _06331_ _06334_ net369 vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ _03289_ net1051 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03115_
+ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__and4_1
XANTENNA__12148__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ net360 net2495 net595 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
X_14587_ net1077 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16326_ clknet_leaf_8_wb_clk_i _02466_ _01134_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13538_ _03093_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09280__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11987__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16257_ clknet_leaf_102_wb_clk_i _02397_ _01065_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13469_ team_02_WB.START_ADDR_VAL_REG\[9\] net1071 net1005 vssd1 vssd1 vccd1 vccd1
+ net223 sky130_fd_sc_hd__a21o_1
XFILLER_0_125_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09568__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15208_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_dready _00021_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.d_ready sky130_fd_sc_hd__dfrtp_1
Xoutput204 net204 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput215 net215 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
X_16188_ clknet_leaf_17_wb_clk_i _02328_ _00996_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10178__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09032__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11288__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ net1157 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_max_cap526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__A1 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _03681_ _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14599__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\] net762 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\]
+ _05214_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a221o_1
XANTENNA__11678__A1 _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ _03584_ _03603_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12611__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\] net811 net911 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a22o_1
XANTENNA__09740__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _05071_ _05074_ _05076_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__nor4_1
XANTENNA__09099__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08513_ net1048 _04202_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09493_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\] net756 net729 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12847__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08444_ _04145_ _04146_ _04147_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__and2_1
XANTENNA__12058__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_A _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1165_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09271__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09559__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__A team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1218_X net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13107__B2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 _05716_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_2
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 _07229_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
XANTENNA__11669__A1 _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 _07225_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12521__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 _07222_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_4
Xfanout464 _07213_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_8
Xfanout475 _07206_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 net489 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_6
XANTENNA__09731__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout497 _06250_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
X_09829_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\] net706 _05344_ _05345_
+ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12919__A1_N _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ _04842_ _06171_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12771_ _06942_ _07039_ _07059_ _07082_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08837__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14510_ net1082 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
X_11722_ net298 net2492 net602 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
X_15490_ clknet_leaf_118_wb_clk_i _01630_ _00298_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14441_ net1214 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
X_11653_ _05336_ _05932_ _05989_ _05380_ _05559_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10604_ _06104_ _06108_ _06120_ _06103_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a211o_1
XANTENNA__09798__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14372_ net1099 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
X_11584_ net395 _06998_ _07070_ _07072_ net384 vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16756__1300 vssd1 vssd1 vccd1 vccd1 _16756__1300/HI net1300 sky130_fd_sc_hd__conb_1
X_16111_ clknet_leaf_41_wb_clk_i _02251_ _00919_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13323_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _03011_ _03010_ net1638
+ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_91_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16042_ clknet_leaf_39_wb_clk_i _02182_ _00850_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13254_ _06415_ _02964_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__or2_1
X_10466_ _04906_ _04908_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_114_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12205_ net359 net2399 net579 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13185_ team_02_WB.instance_to_wrap.top.pc\[4\] net1024 _02944_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01485_ sky130_fd_sc_hd__a22o_1
X_10397_ _05690_ net504 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__and2b_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_209_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12136_ net338 net1813 net469 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12067_ net336 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\] net472 vssd1
+ vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XANTENNA__12431__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09306__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net947 _06523_ _06529_ net606 vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__o211a_4
XFILLER_0_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15826_ clknet_leaf_54_wb_clk_i _01966_ _00634_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15757_ clknet_leaf_40_wb_clk_i _01897_ _00565_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13282__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12969_ team_02_WB.instance_to_wrap.top.pc\[5\] _05695_ vssd1 vssd1 vccd1 vccd1 _07489_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10096__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14708_ net1239 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
X_15688_ clknet_leaf_20_wb_clk_i _01828_ _00496_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ net1224 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14882__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _03840_ net227 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09253__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16309_ clknet_leaf_40_wb_clk_i _02449_ _01117_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _03784_ _03810_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload30 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
Xclkload41 clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_4
XFILLER_0_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload52 clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__inv_12
XFILLER_0_23_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload63 clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__inv_6
XANTENNA__10634__B _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload74 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinv_2
Xclkload85 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_4
Xclkload96 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_167_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09961__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07944_ _03602_ _03605_ _03638_ _03627_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a31o_1
XANTENNA__12341__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07875_ net316 _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09614_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\] net758 net754 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_178_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] net823 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13273__B1 _06618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout638_A _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09476_ _04970_ _04991_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_191_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08427_ _04130_ _04133_ _04128_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_A _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08358_ _04056_ _04064_ _04067_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a31o_2
XFILLER_0_191_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload2 clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__09244__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12516__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ _03966_ _03979_ _03989_ _03970_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_210_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10320_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\] net918 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] net758 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ _05765_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a221o_1
X_10182_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\] net916 net819 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\]
+ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1217 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_4
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_4
Xfanout1237 net1265 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_2
XANTENNA__12251__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14990_ net1154 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
Xfanout250 _06498_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_2
Xfanout1259 net1260 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_4
Xfanout261 _06595_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09704__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 net275 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
Xfanout283 _06657_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
X_13941_ net1164 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
Xfanout294 _06791_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
X_16660_ clknet_leaf_93_wb_clk_i _02779_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13872_ net1165 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
X_15611_ clknet_leaf_33_wb_clk_i _01751_ _00419_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12823_ _04306_ _07340_ _07344_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a21o_1
X_16591_ clknet_leaf_90_wb_clk_i _02710_ _01384_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08684__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15542_ clknet_leaf_49_wb_clk_i _01682_ _00350_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ _05557_ _05604_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09483__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ net240 net2307 net602 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
X_12685_ net273 net2427 net432 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15473_ clknet_leaf_0_wb_clk_i _01613_ _00281_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input91_X net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11636_ net848 _06162_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nand2_1
X_14424_ net1195 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XANTENNA__09235__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11578__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11567_ _05738_ _05911_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__xnor2_1
X_14355_ net1078 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12426__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10250__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ _04569_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13319__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ net1613 net984 net966 _03002_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__a22o_1
X_14286_ net1082 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
Xhold709 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ team_02_WB.instance_to_wrap.top.pc\[8\] net975 _06991_ _04263_ vssd1 vssd1
+ vccd1 vccd1 _06992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ clknet_leaf_124_wb_clk_i _02165_ _00833_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ _02958_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__inv_2
X_10449_ _04630_ _04652_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10002__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ _07009_ net232 _02928_ net976 _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__o221a_1
X_12119_ net269 net2470 net467 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XANTENNA__12161__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ _07519_ _02872_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_127_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07660_ _03380_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__xor2_1
XANTENNA__10856__A2 _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15809_ clknet_leaf_101_wb_clk_i _01949_ _00617_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07591_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__nand2_1
X_16789_ net1333 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_149_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09330_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] net885 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10069__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_192_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09474__A2 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _04714_ _04733_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08212_ _03897_ _03922_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11018__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09192_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] net743 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a221o_1
XANTENNA__09226__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _03852_ _03861_ _03856_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_43_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12336__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09993__X _05510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10241__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _03764_ _03787_ _03791_ _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_141_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13956__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__X _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1128_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 _02624_ vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15267__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ _04326_ _04492_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__or2_4
Xhold25 _02592_ vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_02_WB.instance_to_wrap.ramstore\[13\] vssd1 vssd1 vccd1 vccd1 net1398
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_02_WB.instance_to_wrap.top.a1.data\[7\] vssd1 vssd1 vccd1 vccd1 net1409
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03636_ _03611_ vssd1 vssd1
+ vccd1 vccd1 _03650_ sky130_fd_sc_hd__o21bai_1
Xhold58 team_02_WB.START_ADDR_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_02_WB.instance_to_wrap.ramaddr\[29\] vssd1 vssd1 vccd1 vccd1 net1431
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_208_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout755_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10847__A2 _06344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _03578_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _03507_ _03509_ _03499_ _03501_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout922_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09528_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\] net763 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_158_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09465__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09459_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\] net812 net910 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12470_ net356 net2430 net453 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11421_ net422 _06473_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nand2_1
XANTENNA__12246__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14027__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10232__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ net1201 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
X_11352_ _06104_ _06851_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__nand2_1
XANTENNA__08670__D team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08025__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\] net705 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14071_ net1219 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11283_ _06263_ _06785_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _07540_ _07541_ net230 vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input51_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\] net811 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a221o_1
Xfanout1001 _04263_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_2
Xfanout1012 net1014 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10165_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\] net825 net813 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a22o_1
XANTENNA__10290__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_210_Right_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_2
XANTENNA__16192__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1045 net1046 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
Xfanout1056 team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1056 sky130_fd_sc_hd__buf_2
XFILLER_0_206_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_2
X_14973_ net1161 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
X_10096_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\] net762 net738 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a22o_1
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_4
Xfanout1089 net1094 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_4
XANTENNA_output138_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16712_ net1271 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XANTENNA__10299__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ net1258 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_109_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12929__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16643_ clknet_leaf_95_wb_clk_i _02762_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13855_ net1147 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _07323_ _07324_ _07322_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__mux2_1
X_16574_ clknet_leaf_92_wb_clk_i _00000_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_122_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10998_ _06314_ _06325_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__or2_1
X_13786_ _03276_ _03277_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__nor2_1
XANTENNA__09456__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15525_ clknet_leaf_23_wb_clk_i _01665_ _00333_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12737_ _07260_ _06924_ _07259_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__and3b_1
XANTENNA__09797__Y _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15456_ clknet_leaf_18_wb_clk_i _01596_ _00264_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ net355 net1780 net436 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14407_ net1174 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XANTENNA__12156__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ net948 _07104_ _07106_ net607 vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__o211a_4
XANTENNA__10465__A _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15387_ clknet_leaf_34_wb_clk_i _01527_ _00195_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12599_ net339 net2413 net439 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14338_ net1191 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11995__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14269_ net1204 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
X_16008_ clknet_leaf_20_wb_clk_i _02148_ _00816_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08589__B net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ net1574 net1038 net990 team_02_WB.instance_to_wrap.ramaddr\[1\] vssd1 vssd1
+ vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
Xhold1206 team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1 net2568
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\] net773 net701 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a22o_1
Xhold1217 team_02_WB.instance_to_wrap.top.pad.keyCode\[6\] vssd1 vssd1 vccd1 vccd1
+ net2579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1228 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13476__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _03433_ _03434_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10829__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ net1059 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] net1060 vssd1
+ vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12839__B _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07643_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03334_ _03360_ vssd1 vssd1
+ vccd1 vccd1 _03366_ sky130_fd_sc_hd__or3_1
XANTENNA_wire609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07574_ team_02_WB.instance_to_wrap.top.pad.count\[0\] team_02_WB.instance_to_wrap.top.pad.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__and2b_1
XFILLER_0_165_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09447__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] net739 net715 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_196_Left_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout336_A _06994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\] net824 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\]
+ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a221o_1
XANTENNA__13303__X _03001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09500__Y _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ net971 _04691_ net544 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_153_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12066__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1245_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10214__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _03842_ _03843_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09080__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ _03734_ _03756_ _03736_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_114_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_186_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10517__A1 _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput104 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_168_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] net779 net751 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__A1 _04496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ net356 net1844 net586 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
XANTENNA__09686__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _06302_ _06306_ net368 vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__mux2_1
XANTENNA__13219__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13640_ team_02_WB.instance_to_wrap.top.a1.row2\[15\] _03103_ _03165_ _03117_ team_02_WB.instance_to_wrap.top.a1.row1\[63\]
+ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__a32o_1
X_10852_ _06272_ _06367_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09438__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10783_ _06297_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__or2_1
X_13571_ net1049 _03103_ _03113_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15310_ clknet_leaf_63_wb_clk_i _01453_ _00123_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15141__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09410__Y _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ net293 net2544 net447 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__mux2_1
X_16290_ clknet_leaf_119_wb_clk_i _02430_ _01098_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input99_A wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15241_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[0\]
+ _00054_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12453_ net289 net2098 net451 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__mux2_1
XANTENNA__14980__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10205__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ net424 _06451_ _06900_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__o21ai_2
X_12384_ net271 net1883 net461 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__mux2_1
X_15172_ net1142 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14123_ net1125 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
X_11335_ _06194_ net652 _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _06835_
+ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__a221o_1
XANTENNA__12704__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07594__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14054_ net1212 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
X_11266_ net378 _06539_ _06639_ _06534_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__o22a_1
X_10217_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] net768 net719 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a22o_1
X_13005_ _07460_ _07524_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__and2b_1
XFILLER_0_207_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11197_ _06117_ _06696_ _06699_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__o211ai_1
X_10148_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] net770 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14956_ net1214 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
X_10079_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] net820 net816 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\]
+ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a221o_1
XANTENNA__09677__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13907_ net1167 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XANTENNA__08885__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14887_ net1182 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
X_16626_ clknet_leaf_94_wb_clk_i _02745_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13838_ net1163 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16557_ clknet_leaf_87_wb_clk_i _02681_ _01364_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _03265_ _03266_ net960 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__and3b_1
X_15508_ clknet_leaf_14_wb_clk_i _01648_ _00316_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16488_ clknet_leaf_69_wb_clk_i net1432 _01296_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15439_ clknet_leaf_42_wb_clk_i _01579_ _00247_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14890__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09601__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold325 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12614__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold336 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09048__X _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold358 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold369 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] net910 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout805 _04534_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_4
Xfanout816 _04520_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
X_09862_ _05355_ _05376_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nand2_1
Xfanout827 _04512_ vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
Xfanout838 _04403_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout849 _04186_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
Xhold1003 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net1506 net1038 net990 team_02_WB.instance_to_wrap.ramaddr\[18\] vssd1 vssd1
+ vccd1 vccd1 _02612_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_181_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09793_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\] net764 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a221o_1
Xhold1014 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1047 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _04302_ net931 _04359_ _04368_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__and4_4
XANTENNA__09668__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_163_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _04298_ _04299_ _04300_ _04303_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout453_A _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] _03324_ _03327_ vssd1 vssd1
+ vccd1 vccd1 _03349_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07557_ net1059 vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout718_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10817__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\] net689 net677 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09158_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\] net921 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a22o_1
XANTENNA__09053__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _03824_ _03825_ _03820_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08800__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\] net915 net810 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a221o_1
XANTENNA__12524__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10833__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ net399 _06511_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold870 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11051_ _06151_ _06152_ _06233_ net974 vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__o31a_1
X_10002_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\] net716 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a221o_1
X_14810_ net1096 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_199_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ clknet_leaf_48_wb_clk_i _01930_ _00598_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09659__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1242 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
X_11953_ net289 net2588 net585 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10904_ net975 _06417_ _06418_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and3_1
X_14672_ net1227 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
X_11884_ net278 net2170 net486 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__mux2_1
XANTENNA__08973__A team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16411_ clknet_leaf_85_wb_clk_i _02546_ _01219_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13623_ _03132_ _03172_ _03173_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or4_1
X_10835_ net545 net398 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16342_ clknet_leaf_21_wb_clk_i _02482_ _01150_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13554_ _03107_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09292__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ net1888 net241 net640 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XANTENNA__10977__A1 _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09831__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ net350 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] net556 vssd1
+ vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__mux2_1
X_16273_ clknet_leaf_128_wb_clk_i _02413_ _01081_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13485_ team_02_WB.START_ADDR_VAL_REG\[25\] net1070 net1002 vssd1 vssd1 vccd1 vccd1
+ net209 sky130_fd_sc_hd__a21o_1
X_10697_ _06195_ _06212_ _06213_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ clknet_leaf_104_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[15\]
+ _00037_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_12436_ net361 net1735 net457 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ net1144 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
X_12367_ net330 net2019 net560 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__mux2_1
XANTENNA__12434__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14106_ net1095 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
X_11318_ _06771_ _06818_ net370 vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12298_ net324 net1722 net568 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__mux2_1
X_15086_ net1163 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
X_11249_ _06502_ _06639_ _06752_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_130_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14037_ net1241 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09898__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15988_ clknet_leaf_14_wb_clk_i _02128_ _00796_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08858__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire519_A _05313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14939_ net1085 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14885__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08460_ _04157_ _04162_ _04158_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__o21a_1
XFILLER_0_203_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16609_ clknet_leaf_93_wb_clk_i _02728_ _01402_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08391_ net1593 net1006 net981 _04100_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a22o_1
XANTENNA__12609__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09283__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__Y _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09822__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10129__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ net1058 _04295_ _04297_ net952 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__and4_4
XFILLER_0_115_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09035__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold100 team_02_WB.instance_to_wrap.ramaddr\[28\] vssd1 vssd1 vccd1 vccd1 net1462
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12344__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 _02621_ vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold122 net112 vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 team_02_WB.START_ADDR_VAL_REG\[11\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 net115 vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _02611_ vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_02_WB.START_ADDR_VAL_REG\[30\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 _02618_ vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
X_16736__1282 vssd1 vssd1 vccd1 vccd1 _16736__1282/HI net1282 sky130_fd_sc_hd__conb_1
X_09914_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\] net750 net705 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold199 team_02_WB.instance_to_wrap.top.a1.row1\[107\] vssd1 vssd1 vccd1 vccd1 net1561
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 _07189_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_6
XFILLER_0_186_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout613 net618 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1110_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1208_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout657 net659 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\] net915 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a22o_1
Xfanout668 _05965_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
XANTENNA_fanout570_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_8
X_09776_ net609 _05290_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nand2_1
X_08727_ _04328_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__and2b_1
XANTENNA__08849__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout835_A _04506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14795__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11771__X _07192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08658_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__inv_2
XANTENNA__10120__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07609_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] _03331_ vssd1 vssd1 vccd1
+ vccd1 _03332_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_194_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12519__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ net43 net42 net45 net44 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__or4_1
X_10620_ team_02_WB.instance_to_wrap.top.pc\[29\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _06137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09274__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ net369 _06063_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11081__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10039__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10482_ _05833_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__or2_1
X_13270_ net1634 net982 net964 _02984_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a22o_1
X_12221_ net1824 net277 net612 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
XANTENNA__12254__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11011__X _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ net263 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\] net465 vssd1
+ vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11103_ _06610_ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__or2_1
X_12083_ net1678 net267 net582 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
X_15911_ clknet_leaf_38_wb_clk_i _02051_ _00719_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11034_ net407 _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__nor2_1
XANTENNA__11687__A2 _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_188_Right_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15842_ clknet_leaf_118_wb_clk_i _01982_ _00650_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07591__B team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09176__A_N net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15773_ clknet_leaf_10_wb_clk_i _01913_ _00581_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11439__A2 _06931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ _07484_ _07504_ _07482_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__a21o_1
X_14724_ net1091 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
X_11936_ net354 net1860 net484 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10111__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14655_ net1116 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
X_11867_ net358 net2370 net493 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XANTENNA__12429__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13606_ team_02_WB.instance_to_wrap.top.a1.row1\[19\] _03111_ _03116_ team_02_WB.instance_to_wrap.top.a1.row1\[123\]
+ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a22o_1
X_10818_ _06332_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14586_ net1088 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XANTENNA__09804__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ net345 net2485 net594 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11072__B1 _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16325_ clknet_leaf_29_wb_clk_i _02465_ _01133_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13537_ _03072_ _03078_ _03082_ _03075_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10749_ team_02_WB.instance_to_wrap.top.pc\[22\] team_02_WB.instance_to_wrap.top.pc\[21\]
+ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_41_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16256_ clknet_leaf_17_wb_clk_i _02396_ _01064_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13468_ team_02_WB.START_ADDR_VAL_REG\[8\] _04260_ vssd1 vssd1 vccd1 vccd1 net222
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13281__A1_N _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15207_ clknet_leaf_81_wb_clk_i net1018 _00020_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.i_ready
+ sky130_fd_sc_hd__dfrtp_1
X_12419_ net278 net1831 net454 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XANTENNA__10473__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16187_ clknet_leaf_33_wb_clk_i _02327_ _00995_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12164__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput205 net205 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
X_13399_ team_02_WB.instance_to_wrap.ramload\[28\] net1011 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[28\] sky130_fd_sc_hd__and2_1
Xoutput216 net216 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_11_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15138_ net1157 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
X_15069_ net1253 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
X_07960_ _03656_ _03673_ _03678_ _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_120_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07891_ _03612_ _03613_ _03608_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09630_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\] net903 net887 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a22o_1
XANTENNA__10350__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09561_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\] net830 net896 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\]
+ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a221o_1
X_08512_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\] net979 vssd1 vssd1 vccd1
+ vccd1 _04203_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09492_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] net766 _05000_ _05001_
+ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a2111o_2
XANTENNA__10102__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08443_ _04146_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12339__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout249_A _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ _04072_ _04075_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__xor2_1
XANTENNA__13959__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13311__X _03005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12074__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12563__A0 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08782__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_2
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
Xfanout432 _07229_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_6
Xfanout443 _07225_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_4
Xfanout454 _07221_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_6
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _07213_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
Xfanout476 _07206_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_8
X_09828_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] net782 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a22o_1
Xfanout487 net489 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10341__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12618__A1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] net822 net908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _07112_ _07136_ _07261_ _07271_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__a41o_1
XFILLER_0_96_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09495__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13291__B2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11721_ net310 net2467 net601 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12249__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__A _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14440_ net1112 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11652_ _04482_ _04488_ _04565_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10603_ _04569_ _06110_ net661 _04568_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__a221o_1
XANTENNA__10992__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14371_ net1137 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12773__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11583_ net389 _07071_ net395 vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16110_ clknet_leaf_47_wb_clk_i _02250_ _00918_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input81_A wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ _04174_ _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__or2_1
X_10534_ _06047_ _06050_ net367 vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16041_ clknet_leaf_112_wb_clk_i _02181_ _00849_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11389__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ _04885_ _04905_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nand2_1
X_13253_ net1375 net983 net965 _02972_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11357__A1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ net344 net2213 net578 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ net230 _02941_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a21bo_1
X_10396_ net504 _05690_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2b_1
X_12135_ net331 net1820 net466 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11109__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ net328 net2075 net473 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
X_11017_ net974 _06524_ _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__a211o_1
XANTENNA__10332__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15825_ clknet_leaf_126_wb_clk_i _01965_ _00633_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_15756_ clknet_leaf_126_wb_clk_i _01896_ _00564_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09486__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ _05695_ team_02_WB.instance_to_wrap.top.pc\[5\] vssd1 vssd1 vccd1 vccd1 _07488_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14707_ net1078 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11919_ net290 net1850 net482 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
X_15687_ clknet_leaf_42_wb_clk_i _01827_ _00495_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12159__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12899_ _07372_ _07418_ _07373_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ net1082 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16735__1281 vssd1 vssd1 vccd1 vccd1 _16735__1281/HI net1281 sky130_fd_sc_hd__conb_1
XFILLER_0_172_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11998__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13585__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ net1228 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11596__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16308_ clknet_leaf_14_wb_clk_i _02448_ _01116_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_08090_ _03784_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_122_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16239_ clknet_leaf_41_wb_clk_i _02379_ _01047_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload31 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_max_cap636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload53 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__clkinv_2
Xclkload64 clknet_leaf_88_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_140_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload75 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload75/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload86 clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload86/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload97 clknet_leaf_57_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08764__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12622__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08992_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__and3b_2
XANTENNA_wire541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ _03631_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07874_ _03558_ _03566_ _03589_ _03561_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a22o_2
XANTENNA__10323__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11520__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\] net762 net742 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_178_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09544_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\] net787 _05055_ _05059_
+ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13273__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09475_ net971 _04990_ net543 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12069__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08426_ _04106_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ _04050_ _04051_ _04057_ _04068_ _04044_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__a32oi_1
XANTENNA_fanout700_A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload3 clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08288_ _03962_ _03988_ _03979_ _03970_ _03966_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11339__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] net730 net727 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a221o_1
XANTENNA__09401__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\] net925 net909 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a22o_1
XANTENNA__10841__A _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
Xfanout1216 net1217 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_4
Xfanout1227 net1237 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_2
Xfanout1238 net1240 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_4
Xfanout240 _06282_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1249 net1264 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
Xfanout251 _06498_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_1
Xfanout262 _06595_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_1
XFILLER_0_199_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
X_13940_ net1160 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
Xfanout284 _06766_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_2
XFILLER_0_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout295 _06791_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_1
XANTENNA__09180__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ net1163 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
X_15610_ clknet_leaf_51_wb_clk_i _01750_ _00418_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12822_ _04305_ _07340_ _07344_ team_02_WB.instance_to_wrap.top.a1.state\[2\] vssd1
+ vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22o_1
X_16590_ clknet_leaf_90_wb_clk_i _02709_ _01383_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09468__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ clknet_leaf_40_wb_clk_i _01681_ _00349_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12753_ _05513_ _05904_ _05929_ _07276_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14983__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08029__Y _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11704_ _04291_ net641 _07188_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__or3_4
X_15472_ clknet_leaf_23_wb_clk_i _01612_ _00280_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12684_ net289 net1924 net431 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14423_ net1207 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
X_11635_ _07119_ _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11578__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire630 _05079_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14354_ net1177 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
X_11566_ net376 _06898_ _07055_ _06695_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__a211o_1
XANTENNA__09640__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13305_ team_02_WB.instance_to_wrap.top.pc\[7\] net1054 _07007_ net933 vssd1 vssd1
+ vccd1 vccd1 _03002_ sky130_fd_sc_hd__a22o_1
X_10517_ _04589_ _04608_ _04611_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14285_ net1126 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
X_11497_ _06257_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16024_ clknet_leaf_121_wb_clk_i _02164_ _00832_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13236_ team_02_WB.instance_to_wrap.top.d_ready _03308_ _04268_ _04346_ vssd1 vssd1
+ vccd1 vccd1 _02958_ sky130_fd_sc_hd__or4_1
X_10448_ _04462_ _05963_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12442__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net229 _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nand2_1
X_10379_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\] net808 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12118_ net261 net1940 net467 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13098_ _07464_ _07465_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11591__A1_N net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12049_ net258 net2023 net470 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XANTENNA__10305__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07590_ team_02_WB.instance_to_wrap.top.a1.state\[2\] _03313_ vssd1 vssd1 vccd1 vccd1
+ _03315_ sky130_fd_sc_hd__nand2_1
X_15808_ clknet_leaf_110_wb_clk_i _01948_ _00616_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_16788_ net1332 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_149_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09459__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15739_ clknet_leaf_29_wb_clk_i _01879_ _00547_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ net536 _04775_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08211_ _03922_ _03923_ _03897_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__a21oi_1
X_09191_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] net758 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12617__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11521__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08142_ _03854_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ _03722_ _03763_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12352__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14133__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10661__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11247__B1_N _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] _04330_ net649 team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a22o_1
Xhold15 team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net1377
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 team_02_WB.instance_to_wrap.ramstore\[25\] vssd1 vssd1 vccd1 vccd1 net1388
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_184_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 _02575_ vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03611_ _03637_ vssd1 vssd1
+ vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand3b_1
Xhold48 net181 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_02_WB.instance_to_wrap.top.a1.data\[2\] vssd1 vssd1 vccd1 vccd1 net1421
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ _03545_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_211_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07788_ _03507_ _03509_ _03499_ _03501_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09527_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\] net719 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09458_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\] net832 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\]
+ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09870__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15831__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08409_ _04115_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _04886_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__and2_1
XANTENNA__12527__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _05928_ net660 net657 _05420_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08425__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09622__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11351_ net420 _06348_ _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15981__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08025__B _03746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] net761 net725 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a22o_1
X_14070_ net1106 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11282_ team_02_WB.instance_to_wrap.top.pc\[17\] _06262_ vssd1 vssd1 vccd1 vccd1
+ _06785_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09925__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ _07445_ _07538_ _07539_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__and3_1
XANTENNA__12262__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] net915 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__a22o_1
XANTENNA__15211__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1004 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_2
XANTENNA_input44_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\] net809 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\]
+ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a221o_1
XANTENNA__08041__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
Xfanout1024 net1025 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
Xfanout1046 _04245_ vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_4
X_14972_ net1161 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
X_10095_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] net838 _05609_ _05611_
+ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a211o_1
Xfanout1057 team_02_WB.instance_to_wrap.busy_o vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_2
XANTENNA__09689__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 _00018_ vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1086 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_4
X_16711_ net1270 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
X_13923_ net1234 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XANTENNA__09153__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16642_ clknet_leaf_95_wb_clk_i _02761_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08900__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ net1148 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10289__Y _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _04423_ _07328_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__xor2_1
X_16573_ clknet_leaf_91_wb_clk_i _02697_ _01380_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_13785_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] _03275_
+ net960 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__o21ai_1
X_10997_ net667 _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_122_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15524_ clknet_leaf_35_wb_clk_i _01664_ _00332_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12736_ _06823_ _06851_ _06873_ _06901_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__or4_1
XANTENNA__08915__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15455_ clknet_leaf_62_wb_clk_i _01595_ _00263_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12667_ net359 net1786 net437 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__mux2_1
XANTENNA__12437__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ net1205 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11618_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04347_ net953 _07105_ vssd1
+ vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__a211o_1
XFILLER_0_170_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09613__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15386_ clknet_leaf_53_wb_clk_i _01526_ _00194_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12598_ net330 net2117 net438 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__mux2_1
XANTENNA__12009__Y _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14337_ net1256 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
XANTENNA__11420__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08967__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ net423 _06666_ _07038_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14268_ net1201 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
X_16007_ clknet_leaf_42_wb_clk_i _02147_ _00815_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13219_ net626 net937 net1021 net1398 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12172__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ net1219 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10931__C1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ net847 _04364_ _04370_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__and3_4
Xhold1218 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09144__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ _03302_ net425 _03398_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__a21bo_1
X_08691_ net1059 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04320_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07642_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03360_ _03334_ vssd1 vssd1
+ vccd1 vccd1 _03365_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07573_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] net190 _00017_ vssd1 vssd1
+ vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09312_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\] net759 net752 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\]
+ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09852__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\] net906 vssd1 vssd1
+ vccd1 vccd1 _04760_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12347__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13032__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09174_ _04684_ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08125_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__inv_2
XANTENNA__08958__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1140_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15234__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1238_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A2 _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _03734_ _03756_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout698_A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10391__A _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__C1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput105 wbs_we_i vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_1
XANTENNA_fanout865_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08958_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\] net775 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_205_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09135__A2 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ _03622_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__and2_1
X_08889_ net6 net1029 net986 net2528 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net393 _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__or2_1
XANTENNA__08894__B2 team_02_WB.instance_to_wrap.ramload\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ team_02_WB.instance_to_wrap.top.pc\[30\] _06271_ vssd1 vssd1 vccd1 vccd1
+ _06367_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13570_ net1050 net1051 _03290_ _03103_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__and4b_1
X_10782_ _05534_ net403 vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09843__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12765__B _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ net287 net1738 net446 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__mux2_1
XANTENNA__12257__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15240_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[31\]
+ _00053_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12452_ net278 net1546 net450 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ net424 _06450_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13877__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15171_ net1145 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
X_12383_ net261 net2333 net461 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ net1176 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ net998 _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14053_ net1172 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
X_11265_ _05980_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__xnor2_1
X_13004_ _07461_ _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__nor2_1
XANTENNA__09374__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] net675 _05729_ _05732_
+ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a211o_1
X_11196_ _05041_ net664 _06700_ _06105_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10147_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\] net787 net743 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\]
+ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15877__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14955_ net1123 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10078_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] net922 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13906_ net1153 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
X_14886_ net1212 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
XANTENNA__08885__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10141__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16625_ clknet_leaf_89_wb_clk_i _02744_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13837_ net1155 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16556_ clknet_leaf_91_wb_clk_i _02680_ _01363_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] _03263_
+ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ _06713_ _06741_ _06781_ _07242_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nand4_1
X_15507_ clknet_leaf_51_wb_clk_i _01647_ _00315_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_16487_ clknet_leaf_69_wb_clk_i net1463 _01295_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12167__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] _03221_ vssd1 vssd1 vccd1
+ vccd1 _03222_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15438_ clknet_leaf_48_wb_clk_i _01578_ _00246_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_wire499_A _05828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15369_ clknet_leaf_70_wb_clk_i _01509_ _00182_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[28\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold304 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\] net832 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a22o_1
Xhold359 team_02_WB.instance_to_wrap.ramaddr\[0\] vssd1 vssd1 vccd1 vccd1 net1721
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09365__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 _04534_ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
X_09861_ _05355_ _05376_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__nor2_1
Xfanout817 _04520_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
Xfanout828 _04508_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_8
Xfanout839 _04403_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_0_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08812_ net1558 net1038 net990 team_02_WB.instance_to_wrap.ramaddr\[19\] vssd1 vssd1
+ vccd1 vccd1 _02613_ sky130_fd_sc_hd__a22o_1
XANTENNA__12630__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] net768 net752 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_181_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1004 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1015 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _04302_ _04359_ _04364_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__and3_4
Xhold1048 team_02_WB.instance_to_wrap.ramload\[12\] vssd1 vssd1 vccd1 vccd1 net2410
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1059 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout279_A _06686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ net1063 net1062 _04301_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__and4_1
XFILLER_0_177_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _03324_ _03327_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16032__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1090_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout446_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08628__A1 team_02_WB.START_ADDR_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ team_02_WB.instance_to_wrap.Ren vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_196_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09825__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12077__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout613_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09226_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\] net709 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] net929 net901 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08108_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09088_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\] net865 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13137__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08039_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03744_ _03750_ vssd1 vssd1
+ vccd1 vccd1 _03761_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_92_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold860 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold871 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold893 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net999 _06560_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\] net783 net755 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a22o_1
XANTENNA__10371__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ net1239 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
X_11952_ net279 net2453 net584 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _06136_ _06137_ _06239_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__or3_1
X_14671_ net1199 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
X_11883_ net280 net2149 net488 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16410_ clknet_leaf_105_wb_clk_i _02545_ _01218_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08973__B net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13622_ team_02_WB.instance_to_wrap.top.a1.row1\[3\] _03119_ _03126_ team_02_WB.instance_to_wrap.top.a1.row2\[3\]
+ _03159_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a221o_1
X_10834_ net545 net372 vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09816__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16341_ clknet_leaf_31_wb_clk_i _02481_ _01149_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10765_ net946 _06124_ _06276_ net605 vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__o211a_2
XANTENNA__14991__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12504_ net362 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\] net556 vssd1
+ vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__mux2_1
X_16272_ clknet_leaf_30_wb_clk_i _02412_ _01080_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13484_ team_02_WB.START_ADDR_VAL_REG\[24\] _04260_ vssd1 vssd1 vccd1 vccd1 net208
+ sky130_fd_sc_hd__and2_1
X_10696_ team_02_WB.instance_to_wrap.top.pc\[16\] _06192_ vssd1 vssd1 vccd1 vccd1
+ _06213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15223_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[14\]
+ _00036_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12435_ net344 net1848 net456 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13400__A net2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ net1144 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XANTENNA__09595__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ net334 net2082 net562 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14105_ net1095 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
X_11317_ net521 net406 _06065_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15085_ net1162 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
X_12297_ net320 net1851 net568 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ net1191 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248_ net374 _06503_ _06506_ net379 vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12450__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ net948 _06679_ _06685_ net607 vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__o211a_4
XANTENNA__09325__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15987_ clknet_leaf_56_wb_clk_i _02127_ _00795_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13300__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14938_ net1097 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
XANTENNA__10114__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14869_ net1242 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15062__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16608_ clknet_leaf_96_wb_clk_i _02727_ _01401_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_08390_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__inv_2
XANTENNA__09807__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16539_ clknet_leaf_86_wb_clk_i _02666_ _01346_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09995__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ _04295_ _04297_ net952 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__nand3_4
XANTENNA__12625__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold101 _02622_ vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold112 team_02_WB.instance_to_wrap.top.ru.state\[6\] vssd1 vssd1 vccd1 vccd1 net1474
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _02609_ vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 team_02_WB.instance_to_wrap.ramstore\[11\] vssd1 vssd1 vccd1 vccd1 net1496
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 _02612_ vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 team_02_WB.instance_to_wrap.top.a1.row1\[106\] vssd1 vssd1 vccd1 vccd1 net1518
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold178 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] net729 _05427_ _05429_
+ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__a211o_1
Xfanout603 _07189_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_4
Xhold189 team_02_WB.START_ADDR_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout614 net617 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_6
XANTENNA_fanout396_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09844_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\] net855 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\]
+ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__a221o_1
XANTENNA__12360__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_2
XFILLER_0_95_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10353__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _05965_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_2
X_09775_ net609 _05290_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13980__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ _04344_ _04349_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_197_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10105__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08657_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net997 vssd1 vssd1 vccd1
+ vccd1 _04286_ sky130_fd_sc_hd__nand2b_2
XANTENNA_fanout730_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ _03324_ _03328_ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1
+ vccd1 vccd1 _03331_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_194_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ net104 net71 net105 vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1260_X net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11005__A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10550_ net392 _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] net887 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a22o_1
XANTENNA__12535__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ net390 _05876_ _05995_ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12220_ net2197 net280 net615 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__mux2_1
XANTENNA__09577__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ net266 net1881 net464 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
X_11102_ net417 _06053_ net384 _06101_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__a22o_1
XANTENNA__09329__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ net1931 net260 net580 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
Xhold690 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11136__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net371 _06478_ _06543_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__o21ai_1
X_15910_ clknet_leaf_4_wb_clk_i _02050_ _00718_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12270__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12884__A2 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ clknet_leaf_103_wb_clk_i _01981_ _00649_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14986__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15772_ clknet_leaf_19_wb_clk_i _01912_ _00580_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12984_ _07486_ _07503_ _07485_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08984__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11935_ net361 net1953 net484 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
X_14723_ net1134 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14654_ net1127 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
X_11866_ net342 net2209 net491 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ net1410 net962 _03157_ net1067 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_205_Right_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817_ _05103_ net404 vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08068__A2 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14585_ net1088 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11797_ net338 net2299 net593 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
XANTENNA__13061__A2 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16324_ clknet_leaf_36_wb_clk_i _02464_ _01132_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13536_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] _03061_ _03092_ _03095_
+ net1068 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o221a_1
X_10748_ team_02_WB.instance_to_wrap.top.pc\[20\] _06264_ vssd1 vssd1 vccd1 vccd1
+ _06265_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ clknet_leaf_62_wb_clk_i _02395_ _01063_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13467_ team_02_WB.START_ADDR_VAL_REG\[7\] net1070 net1003 vssd1 vssd1 vccd1 vccd1
+ net221 sky130_fd_sc_hd__a21o_1
X_10679_ net994 _05785_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ clknet_leaf_66_wb_clk_i _01418_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.debounce
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12418_ net280 net2610 net456 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
XANTENNA__09568__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16186_ clknet_leaf_51_wb_clk_i _02326_ _00994_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13398_ net1630 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[27\]
+ sky130_fd_sc_hd__and2_1
Xoutput206 net206 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput217 net217 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ net1157 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12349_ net265 net1809 net561 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ net1251 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ net1136 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12180__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _03575_ _03609_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__xor2_2
XANTENNA_wire531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__C _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10886__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire629_A _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15207__D net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\] net802 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_X clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ team_02_WB.instance_to_wrap.top.a1.data\[6\] net958 vssd1 vssd1 vccd1 vccd1
+ _04202_ sky130_fd_sc_hd__or2_1
XFILLER_0_195_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09491_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] net720 _05005_ _05006_
+ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08700__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ _04135_ _04138_ _04142_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ _04078_ _04080_ _04082_ _04076_ _04075_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__o311a_1
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12355__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout311_A _06840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13975__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
Xfanout411 _05763_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout422 _05715_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout778_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 _07229_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10326__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 _07225_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_6
Xfanout455 _07221_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_4
Xfanout466 net469 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09192__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10877__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout477 _07206_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_4
X_09827_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] net739 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a22o_1
XANTENNA__09731__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\] net903 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08709_ net648 net932 _04337_ _04286_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_87_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09689_ net969 _05205_ _04497_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10839__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11720_ net302 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\] net603 vssd1
+ vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ net665 _07127_ _07136_ _06583_ _07131_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__A2 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10602_ net546 _06117_ _04567_ net658 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09798__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14370_ net1153 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Left_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11582_ _06040_ _06045_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13321_ net1064 _04180_ _04231_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__or3_2
XFILLER_0_91_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10533_ _06048_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nor2_1
XANTENNA__10574__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ clknet_leaf_24_wb_clk_i _02180_ _00848_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13252_ team_02_WB.instance_to_wrap.top.pc\[30\] net1055 _02968_ _02971_ vssd1 vssd1
+ vccd1 vccd1 _02972_ sky130_fd_sc_hd__a22o_1
X_10464_ _04885_ _04905_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__nor2_1
XANTENNA_input74_A wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08044__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12203_ net341 net2086 net577 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13183_ net977 _07397_ _02942_ _07066_ net233 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__o32a_1
X_10395_ _05738_ _05911_ _05736_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a21oi_1
X_12134_ net335 net2379 net467 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12065_ net323 net1803 net470 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
XANTENNA__10317__A0 _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09183__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ _06147_ net653 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] net496
+ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__a221o_1
XANTENNA__09722__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ clknet_leaf_30_wb_clk_i _01964_ _00632_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11817__A0 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15755_ clknet_leaf_17_wb_clk_i _01895_ _00563_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12967_ team_02_WB.instance_to_wrap.top.pc\[6\] _05671_ vssd1 vssd1 vccd1 vccd1 _07487_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13282__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ net276 net1741 net482 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__mux2_1
XANTENNA__10096__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14706_ net1183 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
X_15686_ clknet_leaf_8_wb_clk_i _01826_ _00494_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12898_ _05271_ _06197_ _07417_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ net281 net2232 net492 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
X_14637_ net1121 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11045__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14568_ net1104 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16307_ clknet_leaf_51_wb_clk_i _02447_ _01115_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12175__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ _03074_ _03076_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__or3_1
X_14499_ net1136 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__08461__A2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload10 clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_6
XFILLER_0_70_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload21 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/X sky130_fd_sc_hd__clkbuf_8
X_16238_ clknet_leaf_47_wb_clk_i _02378_ _01046_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload32 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload43 clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_58_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__clkinv_8
Xclkload65 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload65/X sky130_fd_sc_hd__clkbuf_4
Xclkload76 clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload76/X sky130_fd_sc_hd__clkbuf_8
Xclkload87 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__clkinv_4
X_16169_ clknet_leaf_107_wb_clk_i _02309_ _00977_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload98 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__inv_6
XANTENNA__09961__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ net944 _04503_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__and3_4
XFILLER_0_76_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07942_ _03634_ _03637_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nand2_1
X_07873_ _03556_ _03586_ _03587_ _03591_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__o311ai_4
XANTENNA__13019__B _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_wb_clk_i_X clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09612_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\] net710 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\]
+ _05128_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a221o_1
X_09543_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] net771 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_178_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout261_A _06595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13273__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ net970 _04990_ net543 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04119_ _04125_ _04118_ vssd1
+ vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__o31a_1
XANTENNA__12874__A _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1170_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _04055_ _04058_ _04050_ _04051_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_34_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_6
XFILLER_0_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12085__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _03966_ _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_210_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11339__A2 _06830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout895_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\] net827 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1211 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_2
Xfanout1217 net1218 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_2
Xfanout1228 net1230 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_4
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout241 _06282_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_1
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09165__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09704__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout252 _06466_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
Xfanout263 _06595_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout285 _06766_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 _06865_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ net1163 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _03318_ _07342_ _07339_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12752_ _05938_ _05952_ _05958_ _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__or4_1
XANTENNA__10078__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15540_ clknet_leaf_14_wb_clk_i _01680_ _00348_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11275__B2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08039__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11703_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__or3b_2
XFILLER_0_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15471_ clknet_leaf_43_wb_clk_i _01611_ _00279_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12683_ net279 net1855 net430 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__mux2_1
XANTENNA__10856__X _06372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14422_ net1096 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
X_11634_ net654 _07112_ _07120_ net794 vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14353_ net1226 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
Xwire620 _05713_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_2
X_11565_ net393 _06979_ _07054_ net384 vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire631 net632 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15290__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ net1424 net983 net965 _03001_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__a22o_1
X_10516_ _05966_ _06032_ _05967_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21boi_1
X_14284_ net1210 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10250__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11496_ team_02_WB.instance_to_wrap.top.pc\[8\] _06256_ vssd1 vssd1 vccd1 vccd1 _06990_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16023_ clknet_leaf_120_wb_clk_i _02163_ _00831_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13235_ net1053 team_02_WB.instance_to_wrap.top.ru.state\[0\] net982 vssd1 vssd1
+ vccd1 vccd1 _02957_ sky130_fd_sc_hd__o21ba_1
X_10447_ _04462_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__nor2_1
XANTENNA__10002__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09943__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ _07486_ _07503_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__xor2_1
X_10378_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\] net914 _05893_ _05894_
+ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a211o_1
X_12117_ net266 net2162 net468 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
X_13097_ net1027 _02871_ net1025 team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1
+ vccd1 vccd1 _01500_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08996__X _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09156__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ net251 net2175 net471 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__mux2_1
XANTENNA__09604__Y _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15807_ clknet_leaf_59_wb_clk_i _01947_ _00615_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_16787_ net1331 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_205_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13999_ net1220 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12463__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10069__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15738_ clknet_leaf_50_wb_clk_i _01878_ _00546_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15669_ clknet_leaf_40_wb_clk_i _01809_ _00477_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08210_ net2621 net1007 net980 _03927_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11802__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09190_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] net771 _04703_ _04704_
+ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_157_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08141_ _03849_ net227 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload110 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__clkinv_8
X_08072_ _03790_ _03792_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10241__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15783__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12633__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09934__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08412__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap997 _04275_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__buf_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] net789 vssd1 vssd1 vccd1
+ vccd1 _04491_ sky130_fd_sc_hd__or2_2
Xhold16 team_02_WB.instance_to_wrap.ramaddr\[9\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09147__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold27 _02587_ vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03636_ vssd1 vssd1 vccd1
+ vccd1 _03648_ sky130_fd_sc_hd__xnor2_2
Xhold38 team_02_WB.instance_to_wrap.ramstore\[31\] vssd1 vssd1 vccd1 vccd1 net1400
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 net183 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13494__A2 _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _03544_ net329 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07787_ _03507_ _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09526_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] net768 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\] net804 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout810_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout908_A _04524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__A1 _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ _04108_ _04111_ _04102_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ net969 _04904_ _04497_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08339_ _04022_ _04038_ _04027_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_117_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11013__A team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11350_ net375 _06631_ _06849_ net382 vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10232__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\] net737 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12543__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ _06215_ _06216_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_111_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09386__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ _07445_ _07538_ _07539_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10232_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\] net830 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\]
+ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a221o_1
XANTENNA__09925__A2 _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_2
X_10163_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] net899 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__a22o_1
XANTENNA__10940__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1014 _03014_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09138__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 _07348_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
Xfanout1036 _04428_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1047 _04173_ vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input37_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09689__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14971_ net1161 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
X_10094_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\] net766 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\]
+ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__a221o_1
Xfanout1058 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1 vccd1
+ vccd1 net1058 sky130_fd_sc_hd__buf_4
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
X_16710_ net1269 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
X_13922_ net1228 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XANTENNA__10299__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16641_ clknet_leaf_95_wb_clk_i _02760_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13853_ net1150 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12804_ _05835_ _05876_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__xnor2_1
X_16572_ clknet_leaf_87_wb_clk_i _02696_ _01379_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13784_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] _03275_
+ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__and2_1
X_10996_ net422 _06504_ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_122_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15523_ clknet_leaf_9_wb_clk_i _01663_ _00331_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12735_ _06943_ _06963_ _06982_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15454_ clknet_leaf_1_wb_clk_i _01594_ _00262_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12666_ net344 net1688 net435 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14405_ net1117 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
X_11617_ _04263_ net974 team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1 vccd1
+ vccd1 _07105_ sky130_fd_sc_hd__mux2_1
X_12597_ net336 net2548 net441 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__mux2_1
X_15385_ clknet_leaf_124_wb_clk_i _01525_ _00193_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11548_ net423 _06673_ _07038_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14336_ net1102 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12961__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold508 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ net1076 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XANTENNA__12453__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold519 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ team_02_WB.instance_to_wrap.top.pc\[9\] net975 _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\]
+ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__a221o_1
X_13218_ net627 net936 net1020 net1396 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09377__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16006_ clknet_leaf_9_wb_clk_i _02146_ _00814_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09916__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14198_ net1121 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07927__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13149_ net229 _02913_ _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_51_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09129__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1208 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13476__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _03398_ net425 vssd1 vssd1
+ vccd1 vccd1 _03433_ sky130_fd_sc_hd__or3b_1
XANTENNA__11487__B2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__inv_2
XANTENNA__08352__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire611_A _05230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03360_ vssd1 vssd1 vccd1
+ vccd1 _03364_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_205_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07572_ net1064 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] net772 net736 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09301__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12628__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09242_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] net820 net918 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\]
+ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09173_ _04686_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__or3_1
XANTENNA__13125__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08124_ _03778_ _03805_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__nor2_1
XANTENNA__10214__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08055_ _03720_ _03772_ _03773_ _03715_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_189_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12363__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09907__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13164__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10391__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A _07192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\] net735 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_205_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11707__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _03626_ _03629_ _03630_ _03628_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a2bb2o_1
X_08888_ net7 net1033 net989 net1533 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a22o_1
XANTENNA__09540__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ _03521_ _03553_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _06132_ _06240_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719__1351 vssd1 vssd1 vccd1 vccd1 net1351 _16719__1351/LO sky130_fd_sc_hd__conb_1
X_09509_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\] net883 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a22o_1
X_10781_ _05579_ net386 vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12538__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12520_ net273 net1540 net448 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__mux2_1
XANTENNA__11650__A1 _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12451_ net280 net2207 net452 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15211__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11402_ net375 _06691_ _06899_ net380 vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__o22a_1
XANTENNA__11402__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10205__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15170_ net1143 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
X_12382_ net268 net2263 net460 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ net1231 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
X_11333_ team_02_WB.instance_to_wrap.top.pc\[15\] _06261_ vssd1 vssd1 vccd1 vccd1
+ _06834_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12273__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14052_ net1091 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
X_11264_ _05211_ _06016_ _05208_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a21oi_1
X_13003_ _07462_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__nor2_1
X_10215_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\] net788 _05730_ _05731_
+ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a211o_1
XANTENNA__08031__B1 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ _05040_ net658 _06113_ _05038_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08987__A team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\] net758 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10077_ _05587_ _05589_ _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or4_1
X_14954_ net1127 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09531__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ net1254 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
X_14885_ net1175 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
XANTENNA__08885__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload2_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16624_ clknet_leaf_89_wb_clk_i _02743_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13836_ net1154 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XANTENNA__08926__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16555_ clknet_leaf_87_wb_clk_i _02679_ _01362_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_13767_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] _03263_
+ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ _06144_ _06145_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__nor2_1
XANTENNA__12448__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13630__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15506_ clknet_leaf_76_wb_clk_i _01646_ _00314_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11246__B1_N _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _06805_ _06828_ _07241_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_139_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16486_ clknet_leaf_69_wb_clk_i net1473 _01294_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10476__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13698_ net1139 _03220_ _03221_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__nor3_1
XFILLER_0_128_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15437_ clknet_leaf_48_wb_clk_i _01577_ _00245_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12649_ net281 net1863 net436 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15368_ clknet_leaf_70_wb_clk_i _01508_ _00181_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09062__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14319_ net1219 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XANTENNA__12183__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15299_ clknet_leaf_72_wb_clk_i _01443_ _00112_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold327 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14899__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _05356_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__and2_1
Xfanout807 _04534_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_4
XFILLER_0_110_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout818 _04520_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_8
Xfanout829 _04508_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08573__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15821__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ net118 net1038 net990 net1553 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a22o_1
X_09791_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] net731 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a221o_1
Xhold1005 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _04296_ net847 _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__and3_4
Xhold1038 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 team_02_WB.instance_to_wrap.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net2411
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_163_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07624_ _03328_ _03346_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10683__A2 _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12866__B _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ team_02_WB.instance_to_wrap.Wen vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__inv_2
XANTENNA__12358__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout341_A _07030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1083_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\] net749 net705 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_101_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A _06281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09589__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] net835 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09053__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08107_ _03824_ _03825_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__nand2_1
X_09087_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\] net797 _04591_ _04603_
+ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a211o_1
XANTENNA__12093__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08038_ _03744_ _03750_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1
+ vccd1 vccd1 _03760_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold850 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_A _04284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold883 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\] net736 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_110_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09761__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] net919 net899 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11951_ net281 net2566 net586 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _06136_ _06137_ _06239_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__o21ai_1
X_11882_ net271 net2005 net488 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
X_14670_ net1075 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12776__B _06854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10833_ net545 net372 vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13621_ team_02_WB.instance_to_wrap.top.a1.row1\[59\] _03117_ _03123_ team_02_WB.instance_to_wrap.top.a1.row2\[43\]
+ _03158_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12268__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09816__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16340_ clknet_leaf_3_wb_clk_i _02480_ _01148_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13552_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] net1049 vssd1 vssd1 vccd1
+ vccd1 _03107_ sky130_fd_sc_hd__nand2_1
X_10764_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _06278_ _06280_ _04334_
+ team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__o311a_2
XFILLER_0_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09292__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12503_ net356 net1980 net558 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__mux2_1
X_16271_ clknet_leaf_44_wb_clk_i _02411_ _01079_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ team_02_WB.START_ADDR_VAL_REG\[23\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net207 sky130_fd_sc_hd__a21o_1
XFILLER_0_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10695_ _06198_ _06209_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11900__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15222_ clknet_leaf_106_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[13\]
+ _00035_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_12434_ net340 net2405 net454 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09044__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ net1157 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
X_12365_ net326 net1998 net563 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11316_ _05988_ _06816_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__xnor2_1
X_14104_ net1196 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
X_15084_ net1263 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ net313 net1895 net569 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__mux2_1
X_14035_ net1081 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11247_ net422 _06750_ _06355_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__a21boi_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14512__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net998 _06683_ _06684_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__o21ai_1
X_10129_ _05627_ net647 net968 vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__mux2_1
X_15986_ clknet_leaf_55_wb_clk_i _02126_ _00794_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09504__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13300__A1 team_02_WB.instance_to_wrap.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13300__B2 _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14937_ net1090 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XANTENNA__08858__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14868_ net1193 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
X_16607_ clknet_leaf_93_wb_clk_i _02726_ _01400_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_13819_ net1138 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12178__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14799_ net1199 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07818__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16538_ clknet_leaf_87_wb_clk_i _02665_ _01345_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11614__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16469_ clknet_leaf_83_wb_clk_i _02604_ _01277_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
X_09010_ _04295_ _04499_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nand2_1
XANTENNA__11810__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11378__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09035__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold102 net180 vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 team_02_WB.instance_to_wrap.ramstore\[8\] vssd1 vssd1 vccd1 vccd1 net1475
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07597__A2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10050__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 team_02_WB.instance_to_wrap.top.a1.data\[10\] vssd1 vssd1 vccd1 vccd1 net1486
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold135 _02573_ vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 team_02_WB.instance_to_wrap.ramstore\[18\] vssd1 vssd1 vccd1 vccd1 net1508
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 net110 vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09912_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\] net753 net842 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__a221o_1
Xhold179 team_02_WB.instance_to_wrap.top.a1.data\[8\] vssd1 vssd1 vccd1 vccd1 net1541
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12641__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16718__1350 vssd1 vssd1 vccd1 vccd1 net1350 _16718__1350/LO sky130_fd_sc_hd__conb_1
Xfanout604 net606 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_4
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
XANTENNA__09743__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout637 _04454_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_8
X_09843_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\] net891 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__a22o_1
Xfanout648 _04332_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_2
Xfanout659 _06115_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_2
XANTENNA_fanout291_A _06712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _05271_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__and2_1
X_08725_ net648 net932 _04351_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_198_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08849__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _04274_ _04279_ _04280_ net973 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or4_1
XFILLER_0_205_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07607_ _03324_ _03328_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12088__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08587_ _04244_ _04247_ _04248_ net1057 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout723_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_X net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09274__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11720__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ _04718_ _04720_ _04722_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__or4_1
X_10480_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__inv_2
X_09139_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] net730 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12150_ net258 net2032 net462 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
XANTENNA__09982__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ net422 _06069_ net412 vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12551__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12081_ net1667 net251 net582 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
Xhold680 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14332__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold691 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net392 _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or2_1
XANTENNA__09734__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ clknet_leaf_18_wb_clk_i _01980_ _00648_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15771_ clknet_leaf_34_wb_clk_i _01911_ _00579_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13294__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ _03295_ _05671_ _07502_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__o21ai_1
X_14722_ net1129 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
X_11934_ net344 net1707 net484 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
X_14653_ net1206 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
X_11865_ net341 net2068 net491 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ team_02_WB.instance_to_wrap.top.a1.row2\[26\] _03118_ _03150_ _03156_ vssd1
+ vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_107_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10816_ net524 net404 vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11796_ net332 net2434 net592 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
X_14584_ net1195 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16323_ clknet_leaf_25_wb_clk_i _02463_ _01131_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11072__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13535_ _03076_ _03084_ _03093_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__or4_1
XANTENNA__10594__X _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10747_ team_02_WB.instance_to_wrap.top.pc\[19\] team_02_WB.instance_to_wrap.top.pc\[18\]
+ _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10280__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16254_ clknet_leaf_4_wb_clk_i _02394_ _01062_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13466_ team_02_WB.START_ADDR_VAL_REG\[6\] net1070 net1004 vssd1 vssd1 vccd1 vccd1
+ net220 sky130_fd_sc_hd__a21o_1
X_10678_ team_02_WB.instance_to_wrap.top.pc\[15\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _06195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08346__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15205_ clknet_leaf_84_wb_clk_i net1364 _00019_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.flip2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12417_ net270 net2611 net456 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__mux2_1
X_16185_ clknet_leaf_123_wb_clk_i _02325_ _00993_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13397_ net1943 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[26\]
+ sky130_fd_sc_hd__and2_1
Xoutput207 net207 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput218 net218 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_15136_ net1167 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
X_12348_ net257 net2345 net560 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_206_Left_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16022__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12279_ net236 net2144 net568 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__mux2_1
XANTENNA__12461__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15067_ net1250 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09725__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ net1130 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08597__D _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15969_ clknet_leaf_100_wb_clk_i _02109_ _00777_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_08510_ _04201_ net1556 net849 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] net769 net726 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_188_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08441_ _04135_ _04142_ _04138_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13037__B1 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08372_ _04080_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12636__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16405__Q team_02_WB.instance_to_wrap.ramload\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout304_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10023__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12371__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1213_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _05808_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_2
Xfanout412 net415 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09716__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 _05715_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_4
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 _07225_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
Xfanout456 _07221_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_6
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_6
X_09826_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\] net727 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\]
+ _05337_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a221o_1
Xfanout478 net481 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_6
Xfanout489 _07198_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\] net834 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\]
+ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a221o_1
XANTENNA__13276__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16665__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08708_ _04271_ _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09688_ _05198_ _05201_ _05202_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__or4_4
XFILLER_0_179_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09495__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08639_ net1063 net1062 _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__or3_4
XFILLER_0_179_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11650_ _05715_ _06797_ _07134_ _07135_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11581_ net367 _07033_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__nor2_1
XANTENNA__12546__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ _05579_ net403 vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ net1721 net982 net964 _03009_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10262__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10574__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ _05167_ _05168_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and2b_2
X_13251_ _06365_ _02965_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__or2_1
XANTENNA__10014__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12202_ net332 net2191 net577 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
XANTENNA__09955__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13182_ _07388_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__and3_1
X_10394_ _05906_ _05909_ _05783_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__a21bo_1
XANTENNA_input67_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10565__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ net326 net2030 net469 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XANTENNA__12281__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10590__A _05809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09707__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ net317 net2595 net470 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
X_11015_ net999 _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nor2_1
Xfanout990 net993 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_2
X_15823_ clknet_leaf_48_wb_clk_i _01963_ _00631_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_129_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15754_ clknet_leaf_32_wb_clk_i _01894_ _00562_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12966_ team_02_WB.instance_to_wrap.top.pc\[7\] _05627_ vssd1 vssd1 vccd1 vccd1 _07486_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09486__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ net1223 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ net282 net1974 net485 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15685_ clknet_leaf_28_wb_clk_i _01825_ _00493_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12897_ _07374_ _07375_ _07416_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14636_ net1214 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11848_ net270 net1756 net492 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12456__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14567_ net1180 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11779_ net263 net2278 net595 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
XANTENNA__12309__X _07218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ clknet_leaf_77_wb_clk_i _02446_ _01114_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13518_ _03077_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__nor2_1
X_14498_ net1153 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ clknet_leaf_49_wb_clk_i _02377_ _01045_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload11 clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_6
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13449_ _03052_ _03053_ _03041_ _03048_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a2bb2o_1
Xclkload22 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_152_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload33 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload44 clknet_leaf_89_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_58_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10005__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload55 clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__inv_12
XANTENNA__11202__C1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload66 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_6
X_16168_ clknet_leaf_25_wb_clk_i _02308_ _00976_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload77 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_8
XFILLER_0_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload88 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload88/X sky130_fd_sc_hd__clkbuf_4
Xclkload99 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinv_4
X_15119_ net1081 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XANTENNA_max_cap524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12191__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__and3b_2
X_16099_ clknet_leaf_27_wb_clk_i _02239_ _00907_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07941_ _03641_ _03662_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ _03592_ _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08921__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09611_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] net782 net734 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09072__Y _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09542_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] net744 _05044_ _05058_
+ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_178_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ _04980_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nor2_8
XFILLER_0_66_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout254_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08424_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04125_ vssd1 vssd1 vccd1
+ vccd1 _04131_ sky130_fd_sc_hd__nor2_1
XANTENNA__09229__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12874__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _04051_ _04065_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__xor2_2
XFILLER_0_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12366__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1163_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload5 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_22_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ _03962_ _03988_ _03979_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1271_A team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13986__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1207 net1211 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_4
Xfanout1218 net1237 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
Xfanout1229 net1230 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_4
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 _07333_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
Xfanout242 _06282_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 _06466_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_1
Xfanout264 _06595_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_1
Xfanout275 _06740_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08912__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 _06766_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
X_09809_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] net888 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a22o_1
XANTENNA__08912__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 _06865_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_1
XANTENNA__13249__B1 _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12820_ _03318_ _07342_ _07339_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09468__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12751_ _04780_ _05933_ _07272_ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__or4_1
XANTENNA__11275__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15214__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11702_ net2275 net347 net637 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
X_15470_ clknet_leaf_45_wb_clk_i _01610_ _00278_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12682_ net282 net2067 net432 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14421_ net1257 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
X_11633_ net421 _06774_ _07111_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__o21a_1
XANTENNA__12224__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10235__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14352_ net1224 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
X_11564_ net408 _07053_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__or2_1
Xwire632 _05035_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09640__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13303_ team_02_WB.instance_to_wrap.top.pc\[8\] net1054 _06989_ net933 vssd1 vssd1
+ vccd1 vccd1 _03001_ sky130_fd_sc_hd__a22o_1
X_10515_ _04695_ _06031_ net542 _04692_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_190_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11495_ net670 _06976_ _06988_ net672 _06987_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a221o_1
X_14283_ net1125 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
X_16022_ clknet_leaf_22_wb_clk_i _02162_ _00830_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10446_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__nand2_2
X_13234_ team_02_WB.instance_to_wrap.busy_o team_02_WB.instance_to_wrap.top.ru.state\[2\]
+ net1019 _00011_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10377_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] net886 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\]
+ _05885_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a221o_1
X_13165_ _07404_ _07406_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__xnor2_1
X_12116_ net258 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] net466 vssd1
+ vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
X_13096_ _06735_ net234 _02868_ net978 _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_53_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12047_ net255 net1880 net472 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__mux2_1
XANTENNA__12959__B _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15806_ clknet_leaf_4_wb_clk_i _01946_ _00614_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_16786_ net1330 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XANTENNA__09459__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13998_ net1083 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
X_15737_ clknet_leaf_125_wb_clk_i _01877_ _00545_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ team_02_WB.instance_to_wrap.top.pc\[16\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _07469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08131__A2 _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15668_ clknet_leaf_114_wb_clk_i _01808_ _00476_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14619_ net1077 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XANTENNA__12215__A1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__A2 _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ clknet_leaf_41_wb_clk_i _01739_ _00407_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_08140_ net1773 net1007 net980 _03859_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
XANTENNA__10226__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08071_ _03769_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07642__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xclkload100 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__inv_6
Xclkload111 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__09919__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_Left_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11726__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] net790 vssd1 vssd1 vccd1
+ vccd1 _04490_ sky130_fd_sc_hd__nor2_8
Xhold17 _02603_ vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _03615_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__xor2_2
Xhold28 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\] vssd1 vssd1 vccd1 vccd1
+ net1390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14430__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 _02593_ vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13494__A3 _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07855_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] _03575_ _03576_ _03577_ vssd1
+ vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__o211a_1
XANTENNA__09243__B net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_166_Left_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07786_ _03473_ _03497_ _03508_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__inv_2
XFILLER_0_195_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09456_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\] net824 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\]
+ _04972_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09870__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ _04102_ _04108_ _04111_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nand3_1
XANTENNA__12096__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _04897_ _04900_ _04902_ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout803_A _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ _04021_ _04048_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09083__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ _03919_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07633__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_175_Left_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08830__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] net838 _05813_ _05814_
+ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net954 _06782_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\] net876 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a22o_1
X_10162_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] net806 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\]
+ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a221o_1
XANTENNA__15209__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10940__A1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_2
Xfanout1026 net1027 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
X_14970_ net1160 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
X_10093_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] net741 net726 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a22o_1
Xfanout1037 _04428_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_4
Xfanout1048 _04171_ vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_2
XANTENNA__09689__A2 _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 team_02_WB.instance_to_wrap.top.a1.instruction\[13\] vssd1 vssd1 vccd1
+ vccd1 net1059 sky130_fd_sc_hd__buf_2
X_13921_ net1229 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_184_Left_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ clknet_leaf_95_wb_clk_i _02759_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13852_ net1150 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16749__1293 vssd1 vssd1 vccd1 vccd1 _16749__1293/HI net1293 sky130_fd_sc_hd__conb_1
XFILLER_0_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12803_ team_02_WB.instance_to_wrap.top.i_ready net234 vssd1 vssd1 vccd1 vccd1 _07327_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16571_ clknet_leaf_91_wb_clk_i _02695_ _01378_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13783_ _03275_ net960 _03274_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__and3b_1
XANTENNA__12795__A _06102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10995_ net379 _06505_ _06506_ net374 vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11903__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15171__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15522_ clknet_leaf_117_wb_clk_i _01662_ _00330_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12734_ _06284_ _07257_ _06414_ _06035_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07889__A team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453_ clknet_leaf_13_wb_clk_i _01593_ _00261_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12665_ net340 net1729 net435 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10208__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14404_ net1092 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
X_11616_ _07095_ _07096_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09074__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15384_ clknet_leaf_122_wb_clk_i _01524_ _00192_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ net328 net2454 net440 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XANTENNA__10759__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14335_ net1109 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
X_11547_ net377 _06870_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11420__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold509 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09609__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14266_ net1089 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
Xmax_cap228 _03788_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_1
XANTENNA__08513__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ net1000 _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16005_ clknet_leaf_30_wb_clk_i _02145_ _00813_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13217_ _05250_ net936 net1020 net1412 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__a2bb2o_1
X_10429_ _05042_ _05945_ _05038_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14197_ net1241 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_150_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12381__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13148_ _07480_ _07481_ _07508_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_189_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13079_ team_02_WB.instance_to_wrap.top.pc\[22\] net1025 _02856_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01503_ sky130_fd_sc_hd__a22o_1
Xhold1209 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_183_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08888__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07640_ _03332_ _03360_ _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15600__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ net37 net36 net35 net34 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nor4_1
X_16769_ net1313 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_66_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09310_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] net776 _04825_ _04826_
+ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a211o_1
XANTENNA__11813__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09852__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09241_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\] net914 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_90_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09172_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] net818 net943 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\]
+ _04673_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
XANTENNA__09065__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _03778_ _03805_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__nand2_1
XANTENNA__08812__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ _03774_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13164__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1126_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16256__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08956_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\] net699 _04472_ vssd1
+ vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12124__A0 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07907_ _03593_ _03624_ _03594_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__a21o_1
X_08887_ net8 net1029 net986 net2627 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout753_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ _03559_ _03560_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout920_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _03449_ _03477_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09508_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] net833 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ _05024_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _06288_ _06295_ net393 vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__mux2_2
XANTENNA__09843__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09439_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] net773 net729 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a22o_1
XANTENNA__10339__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13232__A1_N net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12450_ net270 net2124 net452 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__inv_2
X_12381_ net260 net1963 net458 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__mux2_1
XANTENNA__12554__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ net1104 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
X_11332_ _04325_ _04354_ _06154_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__a31o_2
XFILLER_0_132_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ net1132 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
X_11263_ net1866 net284 net637 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XANTENNA__12363__A0 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ team_02_WB.instance_to_wrap.top.pc\[19\] _06188_ _07521_ vssd1 vssd1 vccd1
+ vccd1 _07522_ sky130_fd_sc_hd__a21o_1
X_10214_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] net776 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a22o_1
X_11194_ net423 _06693_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10145_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\] net710 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\]
+ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_192_Left_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15623__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14953_ net1218 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
X_10076_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] net805 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\]
+ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__a221o_1
XANTENNA__11510__A2_N net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13904_ net1263 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14884_ net1132 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10141__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16623_ clknet_leaf_89_wb_clk_i _02742_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13835_ net1163 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16554_ clknet_leaf_87_wb_clk_i _02678_ _01361_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_13766_ _03263_ _03264_ net960 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_48_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09295__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13091__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10978_ net953 _06490_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__nand2_1
XANTENNA__09834__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ clknet_leaf_128_wb_clk_i _01645_ _00313_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12717_ _06844_ _06882_ _06895_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__and4_1
X_16485_ clknet_leaf_66_wb_clk_i net1403 _01293_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\]
+ _03217_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15436_ clknet_leaf_3_wb_clk_i _01576_ _00244_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ net269 net2251 net436 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_170_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12464__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15367_ clknet_leaf_72_wb_clk_i _01507_ _00180_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10773__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12579_ net257 net2601 net438 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14318_ net1083 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XANTENNA__11588__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold306 team_02_WB.instance_to_wrap.top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 net1668
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15298_ clknet_leaf_71_wb_clk_i _01442_ _00111_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold317 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold328 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold339 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ net1216 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 _04522_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_8
Xfanout819 _04520_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_2
XANTENNA__11808__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ net1480 net1039 net993 team_02_WB.instance_to_wrap.ramaddr\[21\] vssd1 vssd1
+ vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09790_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] net788 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a22o_1
Xhold1006 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] net931 team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__and3b_2
XPHY_EDGE_ROW_183_Right_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1028 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08672_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] team_02_WB.instance_to_wrap.top.a1.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_163_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07623_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] _03326_ _03330_ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07554_ team_02_WB.instance_to_wrap.top.pc\[6\] vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09286__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09825__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16408__Q team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout334_A _06994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] net769 net753 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_X clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09038__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__B _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09155_ _04656_ _04661_ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__nor3_2
XFILLER_0_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12374__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10199__A2 _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14155__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08106_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09086_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] net822 net814 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\]
+ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08037_ _03741_ _03757_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__xnor2_2
X_16748__1292 vssd1 vssd1 vccd1 vccd1 _16748__1292/HI net1292 sky130_fd_sc_hd__conb_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold840 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11148__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold851 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout870_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _05498_ _05500_ _05502_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or4_1
XANTENNA__10371__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ net1001 net995 _04347_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ net269 net2483 net587 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11320__B2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10901_ net953 _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nand2_1
X_11881_ net264 net2342 net488 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XANTENNA__12549__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ team_02_WB.instance_to_wrap.top.a1.row2\[35\] _03125_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[107\]
+ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a221o_1
X_10832_ net409 _06347_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09816__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13551_ net1049 team_02_WB.instance_to_wrap.top.a1.row2\[12\] _03103_ _03104_ vssd1
+ vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__and4b_1
XFILLER_0_66_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ _04334_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__o21a_1
XANTENNA__15222__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12502_ net358 net2487 net559 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16270_ clknet_leaf_46_wb_clk_i _02410_ _01078_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09029__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input97_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ team_02_WB.START_ADDR_VAL_REG\[22\] _04260_ vssd1 vssd1 vccd1 vccd1 net206
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_101_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10694_ _06195_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15221_ clknet_leaf_106_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[12\]
+ _00034_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_12433_ net332 net2187 net455 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12284__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15152_ net1157 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_12364_ net324 net2217 net560 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14103_ net1208 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
X_11315_ _05295_ _06015_ _05291_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__a21oi_1
X_15083_ net1263 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12295_ net304 net2479 net570 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__mux2_1
X_14034_ net1177 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
X_11246_ _06515_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__o21bai_2
XANTENNA__09201__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ net973 _06681_ _06682_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__a21oi_1
X_10128_ _05629_ _05640_ _05642_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__nor4_2
XFILLER_0_209_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15985_ clknet_leaf_128_wb_clk_i _02125_ _00793_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13300__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\] net709 _05573_ _05575_
+ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a211o_1
X_14936_ net1189 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
XANTENNA__10114__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11311__B2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12967__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_203_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ net1073 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XANTENNA__12459__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16606_ clknet_leaf_95_wb_clk_i _02725_ _01399_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_13818_ net1147 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
XANTENNA__09268__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14798_ net1082 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XANTENNA__09807__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16537_ clknet_leaf_87_wb_clk_i _02664_ _01344_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11614__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13749_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03251_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16468_ clknet_leaf_66_wb_clk_i net1379 _01276_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15419_ clknet_leaf_33_wb_clk_i _01559_ _00227_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12194__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16399_ clknet_leaf_99_wb_clk_i _02534_ _01207_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15669__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09440__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 net151 vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold114 net123 vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 net146 vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold136 net111 vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _02580_ vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _02607_ vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\] net757 net838 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__a22o_1
Xhold169 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12878__A1 _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_186_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09842_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\] net920 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\]
+ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a221o_1
Xfanout638 _04454_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout649 _04332_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_1
XANTENNA__10353__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ net970 net627 net543 vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__o21a_1
XANTENNA__13038__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_A _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _04276_ _04277_ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_198_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10105__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ net1062 _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__nor2_2
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout451_A _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ _03324_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__and2_1
XANTENNA__09259__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__A1 team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08586_ team_02_WB.instance_to_wrap.wb.curr_state\[0\] _04246_ _04243_ vssd1 vssd1
+ vccd1 vccd1 _04248_ sky130_fd_sc_hd__o21a_1
XANTENNA__13055__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12802__A1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08482__A1 _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09207_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\] net818 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09138_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] net743 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08785__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] net739 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11100_ _06607_ _06608_ net418 vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ net1677 net252 net582 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
Xhold670 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _06073_ _06075_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__or2_1
XANTENNA__10344__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15217__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09713__Y _05230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ clknet_leaf_52_wb_clk_i _01910_ _00578_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12982_ _07488_ _07501_ _07487_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13294__B2 _02996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14721_ net1261 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ net340 net2557 net483 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XANTENNA__12279__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14652_ net1192 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
X_11864_ net330 net2398 net490 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
X_13603_ _03132_ _03152_ _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_45_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ net521 net386 _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a21o_1
X_14583_ net1208 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
X_11795_ net336 net2449 net595 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11911__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ clknet_leaf_120_wb_clk_i _02462_ _01130_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13534_ _03072_ _03086_ _03081_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__a21oi_1
X_10746_ team_02_WB.instance_to_wrap.top.pc\[17\] _06262_ vssd1 vssd1 vccd1 vccd1
+ _06263_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16253_ clknet_leaf_4_wb_clk_i _02393_ _01061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ team_02_WB.START_ADDR_VAL_REG\[5\] net1071 net1005 vssd1 vssd1 vccd1 vccd1
+ net219 sky130_fd_sc_hd__a21o_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ net789 _05693_ _06127_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__o22a_2
X_15204_ clknet_leaf_83_wb_clk_i team_02_WB.instance_to_wrap.top.edg2.button_i net1068
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.flip1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ net261 net2466 net456 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16184_ clknet_leaf_122_wb_clk_i _02324_ _00992_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09422__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13396_ net1590 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[25\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__08776__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput208 net208 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
X_15135_ net1167 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ net250 net2059 net561 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
Xoutput219 net219 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__14523__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15066_ net1245 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ net245 net2095 net570 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
X_14017_ net1259 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11229_ team_02_WB.instance_to_wrap.top.pc\[18\] _06263_ team_02_WB.instance_to_wrap.top.pc\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_56_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10335__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09489__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15968_ clknet_leaf_18_wb_clk_i _02108_ _00776_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13285__B2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12189__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ net1181 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
X_15899_ clknet_leaf_30_wb_clk_i _02039_ _00707_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08440_ _04131_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_148_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08371_ _04067_ _04073_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__xor2_2
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11599__A1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09661__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07600__A team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09413__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_wb_clk_i_X clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12652__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1039_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 net404 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
XANTENNA__16421__Q team_02_WB.instance_to_wrap.ramload\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_2
XFILLER_0_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout424 _05715_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1206_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10326__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout435 net437 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_8
Xfanout446 _07224_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_8
Xfanout457 _07221_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\] net735 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a22o_1
XANTENNA__09192__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_8
X_09756_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\] net915 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a22o_1
X_08707_ net1060 _04277_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_1
X_09687_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\] net835 net815 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\]
+ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12099__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A _04506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08638_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04265_ vssd1 vssd1 vccd1
+ vccd1 _04267_ sky130_fd_sc_hd__or2_2
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ _02813_ _04230_ _04180_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_166_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11731__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ _04459_ _06114_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__or2_4
XFILLER_0_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ net2011 net361 net639 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09652__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10531_ _05624_ net385 vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11032__A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ net1717 net983 net965 _02970_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10462_ net525 _05166_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12201_ net334 net2556 net579 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XANTENNA__12562__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _07492_ _07499_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__xor2_1
X_10393_ _05783_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12132_ net321 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\] net466 vssd1
+ vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ net313 net1948 net471 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
X_11014_ _06269_ _06525_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__or2_1
XANTENNA__09183__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12798__A _07321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15174__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 _03320_ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_2
XFILLER_0_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15822_ clknet_leaf_48_wb_clk_i _01962_ _00630_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout991 net993 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ clknet_leaf_113_wb_clk_i _01893_ _00561_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12965_ _05627_ team_02_WB.instance_to_wrap.top.pc\[7\] vssd1 vssd1 vccd1 vccd1 _07485_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14704_ net1225 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
X_11916_ net269 net2555 net485 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ clknet_leaf_35_wb_clk_i _01824_ _00492_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09891__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12896_ _07415_ _07376_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14635_ net1125 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
X_11847_ net263 net1870 net492 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14566_ net1212 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_175_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ net267 net1971 net594 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16305_ clknet_leaf_126_wb_clk_i _02445_ _01113_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13517_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__or4b_2
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10729_ team_02_WB.instance_to_wrap.top.pc\[31\] _06244_ vssd1 vssd1 vccd1 vccd1
+ _06246_ sky130_fd_sc_hd__xor2_1
X_14497_ net1258 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16236_ clknet_leaf_126_wb_clk_i _02376_ _01044_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13448_ _03038_ _02763_ _03051_ _02768_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a31o_1
Xclkload12 clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload23 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_58_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload34 clknet_leaf_110_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_6
Xclkload45 clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__11202__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16167_ clknet_leaf_40_wb_clk_i _02307_ _00975_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12472__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload56 clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_8
XANTENNA__10781__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ team_02_WB.instance_to_wrap.ramload\[8\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[8\] sky130_fd_sc_hd__and2_1
Xclkload67 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_8
Xclkload78 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_6
Xclkload89 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__inv_6
X_15118_ net1080 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XANTENNA__09347__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16098_ clknet_leaf_115_wb_clk_i _02238_ _00906_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15049_ net1235 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
X_07940_ _03645_ _03647_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10308__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_wire634_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _03555_ _03570_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_79_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09610_ _05123_ _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__nand2b_2
XANTENNA__15084__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09541_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] net711 _05056_ _05057_
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09472_ _04982_ _04984_ _04986_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_69_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _04126_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nand2_1
XANTENNA__12647__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout247_A _06372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ _04051_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08285_ _03995_ _03996_ _03974_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or3b_2
Xclkload6 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_6
XFILLER_0_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15237__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1208 net1211 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_2
Xfanout1219 net1223 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
XANTENNA__09544__X _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09165__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 _06282_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_208_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout254 _06466_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11726__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
X_09808_ _05318_ _05320_ _05322_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__or4_1
Xfanout287 _06766_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_1
XANTENNA__10180__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _06865_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\] net743 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\]
+ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12750_ _05123_ _05167_ _05207_ _07273_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11701_ net607 _07184_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__and3_2
XANTENNA__10483__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12681_ net270 net2471 net433 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__mux2_1
XANTENNA__12557__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14420_ net1238 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
XANTENNA__13242__A _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11632_ net665 net378 _06534_ _07116_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__o311a_1
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09625__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ net1219 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ _07015_ _07052_ net367 vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire611 _05230_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15230__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire622 _05689_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_2
Xwire633 _04860_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_1
X_13302_ net1378 net985 net966 _03000_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__a22o_1
X_10514_ _05968_ _06030_ _05969_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__a21o_1
Xwire644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_2
X_14282_ net1188 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
X_11494_ _05559_ _05924_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__xnor2_1
X_16021_ clknet_leaf_22_wb_clk_i _02161_ _00829_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15169__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ net1057 team_02_WB.instance_to_wrap.top.ru.state\[4\] net1372 vssd1 vssd1
+ vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ net837 _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__nor2_1
XANTENNA__12292__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13164_ team_02_WB.instance_to_wrap.top.pc\[8\] net1023 _02927_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01489_ sky130_fd_sc_hd__a22o_1
X_10376_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\] net828 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12115_ net251 net2332 net468 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
X_13095_ net231 _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_53_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ net236 net2060 net473 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XANTENNA__11499__B1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10171__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15805_ clknet_leaf_12_wb_clk_i _01945_ _00613_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_16785_ net1329 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_205_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13997_ net1121 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09901__Y _05418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15736_ clknet_leaf_121_wb_clk_i _01876_ _00544_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12948_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10474__A1 _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15667_ clknet_leaf_47_wb_clk_i _01807_ _00475_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12467__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ net505 _05671_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14618_ net1088 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
X_15598_ clknet_leaf_44_wb_clk_i _01738_ _00406_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14549_ net1242 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08070_ _03765_ _03787_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__nor2_2
Xclkload101 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_12
Xclkload112 clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__inv_6
XFILLER_0_126_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16219_ clknet_leaf_32_wb_clk_i _02359_ _01027_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15079__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08972_ _04482_ _04488_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__nor2_2
X_07923_ _03618_ _03637_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__and2_1
XANTENNA__09147__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1
+ net1380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 team_02_WB.instance_to_wrap.top.a1.data\[6\] vssd1 vssd1 vccd1 vccd1 net1391
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07854_ _03304_ _03568_ _03543_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a21o_1
XANTENNA__10162__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ _03471_ net366 _03472_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout364_A _07107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ _05038_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_84_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09855__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12885__B _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09455_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\] net926 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a22o_1
XANTENNA__12377__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08406_ _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] net912 net901 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\]
+ _04888_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08337_ _04046_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2_1
XANTENNA__11414__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08268_ _03945_ _03948_ _03957_ _03960_ _03935_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a41o_1
XFILLER_0_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout998_A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ _03910_ _03867_ _03905_ _03913_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_197_Right_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09386__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10230_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\] net818 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\] net903 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a22o_1
XANTENNA__14621__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1005 _04259_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_2
XANTENNA__09138__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1027 _07338_ vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_4
X_10092_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] net721 net843 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_2
X_13920_ net1234 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13851_ net1138 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15225__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12802_ _04264_ net551 _07232_ _07235_ _07325_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__a2111oi_2
X_13782_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ _03271_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and3_1
X_16570_ clknet_leaf_87_wb_clk_i _02694_ _01377_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ _06310_ _06335_ net393 vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__mux2_1
XANTENNA__09846__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12733_ _06427_ _06603_ _07256_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__or3_1
XANTENNA__09310__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15521_ clknet_leaf_102_wb_clk_i _01661_ _00329_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12287__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15452_ clknet_leaf_19_wb_clk_i _01592_ _00260_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12664_ net333 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] net434 vssd1
+ vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14403_ net1132 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11615_ net668 _07098_ _07099_ net665 _07102_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10883__X _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15383_ clknet_leaf_115_wb_clk_i _01523_ _00191_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_154_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12595_ net324 net1730 net438 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14334_ net1188 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
X_11546_ net396 _06960_ _07036_ net383 vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08821__B2 team_02_WB.instance_to_wrap.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13158__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14265_ net1099 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11477_ team_02_WB.instance_to_wrap.top.pc\[9\] _06257_ vssd1 vssd1 vccd1 vccd1 _06972_
+ sky130_fd_sc_hd__xnor2_1
X_16004_ clknet_leaf_36_wb_clk_i _02144_ _00812_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13216_ net1571 net1021 net939 _05205_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a22o_1
X_10428_ _05082_ _05944_ _05081_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09377__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14196_ net1239 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ _07480_ _07481_ _07508_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__or3_1
X_10359_ _05869_ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__nor2_8
XFILLER_0_21_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09129__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ net978 _07429_ _02854_ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__o31ai_1
XANTENNA__11366__S net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ net312 net1769 net475 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux2_1
XANTENNA__08888__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11892__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__and2_1
X_16768_ net1312 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09301__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ clknet_leaf_40_wb_clk_i _01859_ _00527_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12197__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16699_ net1266 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_201_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09240_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\] net832 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_X clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09171_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\] net827 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\]
+ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08122_ _03815_ _03816_ _03801_ _03803_ _03807_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08475__A_N team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ _03731_ _03768_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__Y _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11175__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__Y _04339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] net706 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_A _07204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout579_A _07214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_205_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _03596_ _03597_ _03624_ _03587_ _03586_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__a2111o_1
X_08886_ net9 net1029 net986 net2477 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__o22a_1
XANTENNA__08879__B2 net2514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09540__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ _03525_ _03534_ _03527_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_98_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout746_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07768_ _03442_ _03486_ _03487_ _03440_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a22o_1
XANTENNA__09828__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\] net893 net873 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout913_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ _03392_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_121_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09438_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\] net741 _04953_ _04954_
+ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13214__A2_N net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ _06794_ _06897_ net397 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_97_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12380_ net248 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\] net459 vssd1
+ vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11331_ _04325_ _06161_ _06248_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__and3b_1
XANTENNA__09359__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14050_ net1130 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_11262_ net948 _06759_ _06765_ net607 vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_37_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13001_ _07463_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__and2b_1
X_10213_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\] net707 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12570__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _06037_ _06698_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_X clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10374__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__Y _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\] net726 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13312__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\] net829 net899 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__a22o_1
X_14952_ net1110 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XANTENNA__10126__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ net1254 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
X_14883_ net1132 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
XANTENNA__11914__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16622_ clknet_leaf_97_wb_clk_i _02741_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13834_ net1162 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13765_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03264_ sky130_fd_sc_hd__a21o_1
X_16553_ clknet_leaf_90_wb_clk_i _02677_ _01360_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_10977_ _06122_ _06482_ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_48_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13091__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ clknet_leaf_23_wb_clk_i _01644_ _00312_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12716_ _06929_ _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__nor2_1
X_13696_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] _03217_ net1604 vssd1 vssd1
+ vccd1 vccd1 _03220_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16484_ clknet_leaf_71_wb_clk_i net1477 _01292_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12647_ net263 net2069 net436 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15435_ clknet_leaf_113_wb_clk_i _01575_ _00243_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ clknet_leaf_72_wb_clk_i _01506_ _00179_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[25\]
+ sky130_fd_sc_hd__dfstp_2
X_12578_ net250 net1598 net440 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11529_ _05649_ _06110_ net660 _05647_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__a221o_1
X_14317_ net1120 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15297_ clknet_leaf_70_wb_clk_i _01441_ _00110_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold307 team_02_WB.instance_to_wrap.top.a1.row1\[1\] vssd1 vssd1 vccd1 vccd1 net1669
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 team_02_WB.instance_to_wrap.top.a1.row1\[105\] vssd1 vssd1 vccd1 vccd1 net1680
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net1111 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
Xhold329 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_185_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ net1132 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XANTENNA__12480__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 _04522_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_2
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire547_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16769__1313 vssd1 vssd1 vccd1 vccd1 _16769__1313/HI net1313 sky130_fd_sc_hd__conb_1
XANTENNA__09770__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ _04302_ net931 net847 _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__and4_4
Xhold1007 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08671_ net1058 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__and4_1
XANTENNA__11824__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710__1269 vssd1 vssd1 vccd1 vccd1 _16710__1269/HI net1269 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_163_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15092__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__or2_2
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07603__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__A0 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07553_ team_02_WB.instance_to_wrap.top.pc\[12\] vssd1 vssd1 vccd1 vccd1 _03294_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_200_Right_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09223_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\] net681 net838 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12655__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] net704 _04662_ _04663_
+ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09589__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08105_ _03796_ _03821_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09085_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\] net880 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_15_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1236_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ _03741_ _03743_ _03751_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or3_2
Xinput90 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
Xhold830 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold841 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout696_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12390__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12243__X _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1024_X net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold896 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] net927 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout863_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ _04268_ _04346_ _04283_ net998 vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08869_ net1057 team_02_WB.instance_to_wrap.wb.prev_BUSY_O net1031 vssd1 vssd1 vccd1
+ vccd1 _04431_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net837 _06376_ _06414_ net669 _06412_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o221a_2
XANTENNA__11734__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ net267 net2248 net487 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ net398 _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nand2_1
XANTENNA__11608__B1 _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] net1049 vssd1 vssd1 vccd1
+ vccd1 _03105_ sky130_fd_sc_hd__nor2_1
X_10762_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04334_ vssd1 vssd1 vccd1
+ vccd1 _06279_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12501_ net345 net1999 net558 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__mux2_1
X_13481_ team_02_WB.START_ADDR_VAL_REG\[21\] net1070 net1002 vssd1 vssd1 vccd1 vccd1
+ net205 sky130_fd_sc_hd__a21o_1
XANTENNA__10874__A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10693_ team_02_WB.instance_to_wrap.top.pc\[15\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _06210_ sky130_fd_sc_hd__or2_1
X_15220_ clknet_leaf_98_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[11\]
+ _00033_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_12432_ net336 net2268 net457 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_33_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15151_ net1159 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12363_ net320 net2364 net560 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14102_ net1107 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11314_ net1658 net301 net639 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
X_15082_ net1254 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
X_12294_ net297 net2016 net571 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14033_ net1231 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
XANTENNA__11909__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ net413 _06513_ _06748_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__o21ba_1
XANTENNA__15177__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10347__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09752__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ team_02_WB.instance_to_wrap.top.pc\[21\] _06265_ vssd1 vssd1 vccd1 vccd1
+ _06683_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08960__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\] net832 net897 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\]
+ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_42_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15984_ clknet_leaf_23_wb_clk_i _02124_ _00792_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_180_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09903__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14935_ net1185 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
X_10058_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\] net761 _05560_ _05574_
+ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a211o_1
XFILLER_0_203_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14866_ net1185 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16605_ clknet_leaf_95_wb_clk_i _02724_ _01398_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_13817_ net1138 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
XANTENNA__16509__Q team_02_WB.START_ADDR_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14797_ net1126 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_34_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16536_ clknet_leaf_86_wb_clk_i _02663_ _01343_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13748_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03251_ net950 vssd1
+ vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_46_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10784__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12475__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16467_ clknet_leaf_69_wb_clk_i net1425 _01275_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\] _03198_ vssd1 vssd1 vccd1
+ vccd1 _03210_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13293__A1_N _06883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15418_ clknet_leaf_53_wb_clk_i _01558_ _00226_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16398_ clknet_leaf_88_wb_clk_i _02533_ _01206_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11378__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ clknet_leaf_74_wb_clk_i _01489_ _00162_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__15270__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold104 _02582_ vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16396__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold115 _02619_ vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _02578_ vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09991__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold137 _02608_ vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11819__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__B1 _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold148 net120 vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\] net765 net737 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a22o_1
Xhold159 team_02_WB.START_ADDR_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 _06281_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_2
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] net927 net924 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a22o_1
XANTENNA__09743__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 net640 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkload14_A clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _05274_ _05284_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__nor4_2
X_08723_ team_02_WB.instance_to_wrap.top.a1.instruction\[5\] _04266_ _04289_ _04346_
+ _04269_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_198_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08654_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ _04262_ team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ _04283_ sky130_fd_sc_hd__or4bb_4
X_07605_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03325_ _03322_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1 vccd1 _03328_
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__09259__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ net1 _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout444_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1186_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12385__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] net908 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09137_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\] net747 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1141_X net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09068_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\] net727 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\]
+ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a221o_1
XANTENNA__09982__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08019_ _03740_ _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nor2_1
XANTENNA__11729__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10329__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11526__C1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold671 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11030_ net384 _06537_ _06538_ _06540_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__a31o_1
Xhold682 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A2 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ _07490_ _07500_ _07489_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13294__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14720_ net1105 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13245__A _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ net333 net2042 net483 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
X_11863_ net335 net1757 net493 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
X_14651_ net1077 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_200_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15233__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814_ _05231_ net386 vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
X_13602_ team_02_WB.instance_to_wrap.top.a1.row1\[2\] _03119_ _03122_ team_02_WB.instance_to_wrap.top.a1.row2\[10\]
+ _03149_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_45_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ net1107 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
X_11794_ net325 net2498 net593 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16321_ clknet_leaf_104_wb_clk_i _02461_ _01129_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12295__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13533_ _03075_ _03077_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__nor2_1
X_10745_ team_02_WB.instance_to_wrap.top.pc\[16\] team_02_WB.instance_to_wrap.top.pc\[15\]
+ _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__and3_1
X_16768__1312 vssd1 vssd1 vccd1 vccd1 _16768__1312/HI net1312 sky130_fd_sc_hd__conb_1
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14076__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10280__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ team_02_WB.START_ADDR_VAL_REG\[4\] _04260_ vssd1 vssd1 vccd1 vccd1 net218
+ sky130_fd_sc_hd__and2_1
X_16252_ clknet_leaf_21_wb_clk_i _02392_ _01060_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ net994 _05740_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12415_ net265 net2293 net456 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
X_15203_ net1250 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16183_ clknet_leaf_115_wb_clk_i _02323_ _00991_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13395_ net1696 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[24\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__14804__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12346_ net254 net1706 net562 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__mux2_1
X_15134_ net1165 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
Xoutput209 net209 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_116_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15065_ net1166 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
X_12277_ net240 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] net571 vssd1
+ vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__mux2_1
X_14016_ net1105 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XANTENNA__09186__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _06221_ _06222_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16724__1279 vssd1 vssd1 vccd1 vccd1 _16724__1279/HI net1279 sky130_fd_sc_hd__conb_1
X_11159_ _06405_ _06665_ net413 vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15967_ clknet_leaf_62_wb_clk_i _02107_ _00775_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10099__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14918_ net1218 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ clknet_leaf_19_wb_clk_i _02038_ _00706_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14849_ net1260 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
X_08370_ _04073_ _04079_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09110__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16519_ clknet_leaf_127_wb_clk_i _02653_ _01326_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07600__B team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10023__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09964__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__A _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09716__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 net404 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout425 _03427_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_2
XANTENNA_fanout394_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_8
Xfanout447 _07224_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_4
X_09824_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\] net758 _05340_ vssd1
+ vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a21o_1
Xfanout458 _07220_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1101_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout469 _07211_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_4
XANTENNA__12888__B _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09755_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\] net895 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout561_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ _04308_ _04330_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__or2_1
XANTENNA__11287__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] net909 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04265_ vssd1 vssd1 vccd1
+ vccd1 _04266_ sky130_fd_sc_hd__nor2_2
XFILLER_0_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout826_A _04512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07998__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ net2630 _04235_ _04225_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XANTENNA__09101__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08499_ team_02_WB.instance_to_wrap.top.a1.data\[9\] net958 _04193_ vssd1 vssd1 vccd1
+ vccd1 _04194_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10530_ _06045_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_118_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10262__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10461_ net525 _05166_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12200_ net327 net2185 net577 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
XANTENNA__10014__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13180_ net1026 _02940_ net1023 team_02_WB.instance_to_wrap.top.pc\[5\] vssd1 vssd1
+ vccd1 vccd1 _01486_ sky130_fd_sc_hd__a2bb2o_1
X_10392_ net412 net608 vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__nand2_1
XANTENNA__11463__A2_N net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net318 net2570 net466 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09168__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net305 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\] net472 vssd1
+ vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XANTENNA__09707__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15228__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A2 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ team_02_WB.instance_to_wrap.top.pc\[26\] _06268_ vssd1 vssd1 vccd1 vccd1
+ _06525_ sky130_fd_sc_hd__nor2_1
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_4
X_15821_ clknet_leaf_48_wb_clk_i _01961_ _00629_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout981 _03320_ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__buf_2
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15752_ clknet_leaf_24_wb_clk_i _01892_ _00560_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12964_ _07482_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__nor2_1
XANTENNA__09340__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1190 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
X_14703_ net1197 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
X_11915_ net264 net2546 net485 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ clknet_leaf_27_wb_clk_i _01823_ _00491_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _07377_ _07380_ _07413_ _06205_ _05356_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_200_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11922__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15190__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14634_ net1178 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
X_11846_ net266 net1933 net492 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ net257 net2216 net592 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
X_14565_ net1172 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16304_ clknet_leaf_23_wb_clk_i _02444_ _01112_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13516_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__or4b_2
X_10728_ _06244_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__inv_2
XANTENNA__10253__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07926__A_N team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14496_ net1102 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16235_ clknet_leaf_14_wb_clk_i _02375_ _01043_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13447_ _03038_ _02763_ _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a21oi_1
X_10659_ net994 _05442_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nand2_1
XANTENNA__14534__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload13 clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/X sky130_fd_sc_hd__clkbuf_8
Xclkload24 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_8
XFILLER_0_180_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload35 clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_8
XANTENNA__10005__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_58_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13378_ team_02_WB.instance_to_wrap.ramload\[7\] net1014 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[7\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11202__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16166_ clknet_leaf_8_wb_clk_i _02306_ _00974_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload57 clknet_leaf_81_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_16
Xclkload68 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_8
Xclkload79 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinv_8
X_15117_ net1074 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XANTENNA_max_cap624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12329_ net312 net2594 net566 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
X_16097_ clknet_leaf_103_wb_clk_i _02237_ _00905_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09159__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15048_ net1246 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07870_ _03554_ _03570_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__nand2_1
XANTENNA_wire627_A _05289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09540_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\] net783 net752 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_183_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09331__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09471_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\] net918 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ _04121_ _04125_ _04114_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12769__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__Y _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _04046_ _04049_ _04058_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_178_Right_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08284_ _03974_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__xnor2_1
Xclkload7 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12663__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13194__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout776_A _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1211 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_4
Xfanout233 net235 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 net247 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 _06466_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlymetal6s2s_1
X_16767__1311 vssd1 vssd1 vccd1 vccd1 _16767__1311/HI net1311 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_208_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09570__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 net268 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
X_09807_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\] net827 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a221o_1
Xfanout277 net279 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
Xfanout288 net291 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout943_A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ _03305_ _03703_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 _06865_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_1
XANTENNA__13249__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\] net746 net739 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a22o_1
XANTENNA__09322__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ _05180_ _05182_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor4_1
XANTENNA__08381__A_N team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14619__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11742__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11700_ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] _04347_ net953 _07185_ vssd1
+ vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__a211o_1
X_12680_ net263 net1923 net433 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__mux2_1
XANTENNA__11680__A1 _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10483__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11631_ net670 _07117_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11562_ _06290_ _06292_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_7_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14350_ net1075 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16723__1278 vssd1 vssd1 vccd1 vccd1 _16723__1278/HI net1278 sky130_fd_sc_hd__conb_1
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire623 _05463_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_2
X_10513_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__inv_2
Xwire634 _04732_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_2
X_13301_ team_02_WB.instance_to_wrap.top.pc\[9\] net1054 _06970_ net933 vssd1 vssd1
+ vccd1 vccd1 _03000_ sky130_fd_sc_hd__a22o_1
X_14281_ net1231 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
X_11493_ _06985_ _06986_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__nand2_1
Xwire645 _05898_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_21_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16020_ clknet_leaf_3_wb_clk_i _02160_ _00828_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13232_ net644 net938 net1019 net1654 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a2bb2o_1
X_10444_ _04569_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__xor2_1
XANTENNA_input72_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13185__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13077__A1_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ net229 _02926_ _02925_ _02923_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a211o_1
X_10375_ _05887_ _05888_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12114_ net253 net2081 net467 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
X_16746__1291 vssd1 vssd1 vccd1 vccd1 _16746__1291/HI net1291 sky130_fd_sc_hd__conb_1
X_13094_ _07463_ _07520_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11917__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11499__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12045_ net244 net2625 net471 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
XANTENNA__09454__Y _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15804_ clknet_leaf_20_wb_clk_i _01944_ _00612_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_16784_ net1328 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
X_13996_ net1215 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XANTENNA__13645__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ clknet_leaf_119_wb_clk_i _01875_ _00543_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12947_ team_02_WB.instance_to_wrap.top.pc\[16\] _06194_ vssd1 vssd1 vccd1 vccd1
+ _07467_ sky130_fd_sc_hd__nand2_1
XANTENNA__14529__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13660__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11505__X _06998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15666_ clknet_leaf_52_wb_clk_i _01806_ _00474_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12878_ _05695_ net500 _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_158_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ net1091 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
X_11829_ net334 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\] net589 vssd1
+ vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
X_15597_ clknet_leaf_49_wb_clk_i _01737_ _00405_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07627__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10226__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14548_ net1241 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12483__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14479_ net1221 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XANTENNA__10792__A _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload102 clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__inv_8
Xclkload113 clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload113/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__07577__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16218_ clknet_leaf_53_wb_clk_i _02358_ _01026_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09919__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_188_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16149_ clknet_leaf_31_wb_clk_i _02289_ _00957_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15824__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] net754 _04483_ _04485_
+ _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15095__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ _03639_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__or2_1
Xhold19 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net1381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _03304_ _03543_ net329 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__nand3_1
X_07784_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] _03506_ _03504_ _03503_ vssd1
+ vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09523_ _05016_ _05036_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12658__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_203_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14439__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A _07087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1099_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08405_ _04090_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09385_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\] net810 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\]
+ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10217__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _04019_ _04038_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11414__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ _03963_ _03982_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__or2_1
XANTENNA__12393__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ _03909_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__nor2_1
XANTENNA__12914__A1 _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09791__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\] net883 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\]
+ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1008 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1017 team_02_WB.instance_to_wrap.top.ru.next_iready vssd1 vssd1 vccd1 vccd1
+ net1017 sky130_fd_sc_hd__clkbuf_2
X_10091_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\] net781 _05606_ _05607_
+ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a211o_1
Xfanout1028 _07337_ vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_4
Xfanout1039 net1046 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09543__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13850_ net1148 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _07324_ _07323_ _07322_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__mux2_1
X_13781_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\]
+ _03269_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\] vssd1
+ vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a31o_1
XANTENNA__12568__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ _06328_ _06341_ net408 vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11102__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14349__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15520_ clknet_leaf_18_wb_clk_i _01660_ _00328_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12732_ _06485_ _07255_ _06647_ _06660_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_26_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15451_ clknet_leaf_33_wb_clk_i _01591_ _00259_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12663_ net337 net2593 net436 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402_ net1129 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_172_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _05832_ net663 _07100_ net836 _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__o221a_1
XANTENNA__10208__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ clknet_leaf_0_wb_clk_i _01522_ _00190_ vssd1 vssd1 vccd1 vccd1 team_02_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09074__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ net318 net2511 net438 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__mux2_1
XANTENNA__08634__X _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ net1181 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ net396 _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14264_ net1196 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11476_ net946 _06970_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__or2_1
XANTENNA__11169__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16003_ clknet_leaf_26_wb_clk_i _02143_ _00811_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13215_ net1434 net1022 net939 _05164_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a22o_1
X_10427_ _05127_ _05943_ _05123_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__o21ba_1
X_14195_ net1080 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XANTENNA__09782__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\] net677 _05871_ _05873_
+ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13146_ team_02_WB.instance_to_wrap.top.pc\[11\] net1025 _02912_ vssd1 vssd1 vccd1
+ vccd1 _01492_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ net231 _02853_ _06653_ net234 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__o2bb2a_1
X_10289_ _05795_ _05800_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__nor3_2
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09534__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ net305 net1826 net477 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08888__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12986__B _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16767_ net1311 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__12478__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ net1082 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11235__X _06740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15718_ clknet_leaf_7_wb_clk_i _01858_ _00526_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ net138 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_157_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15649_ clknet_leaf_101_wb_clk_i _01789_ _00457_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] net916 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09065__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08121_ _03815_ _03816_ _03801_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16766__1310 vssd1 vssd1 vccd1 vccd1 _16766__1310/HI net1310 sky130_fd_sc_hd__conb_1
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08704__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ _03718_ _03772_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09773__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13338__A net2397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\] net787 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ net316 _03597_ _03626_ _03587_ _03586_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_90_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13057__B _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ net10 net1033 net989 net1552 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout474_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16722__1277 vssd1 vssd1 vccd1 vccd1 _16722__1277/HI net1277 sky130_fd_sc_hd__conb_1
X_07836_ _03525_ _03527_ _03535_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_108_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13085__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _03474_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout739_A _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\] net914 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__a221o_1
X_07698_ _03378_ _03387_ _03395_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745__1290 vssd1 vssd1 vccd1 vccd1 _16745__1290/HI net1290 sky130_fd_sc_hd__conb_1
X_09437_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] net749 net701 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_A _04524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_X net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09368_ _04878_ _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nor2_2
XANTENNA__09056__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ _04006_ _04029_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] net830 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a221o_1
XANTENNA__10071__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11330_ _06198_ _06209_ _06211_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ _04284_ _06760_ _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_37_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10212_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\] net740 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__a22o_1
X_13000_ _07464_ _07519_ _07465_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__o21bai_2
XANTENNA__09764__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _06432_ _06639_ _06697_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11571__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\] net718 _05652_ _05653_
+ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13248__A _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09516__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__B2 _03005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\] net812 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\]
+ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a221o_1
XANTENNA_input35_A gpio_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ net1180 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XANTENNA__15236__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ net1253 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10677__A2 _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14882_ net1153 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
X_16621_ clknet_leaf_97_wb_clk_i _02740_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13833_ net1162 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
XANTENNA__12298__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16552_ clknet_leaf_87_wb_clk_i _02676_ _01359_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[111\]
+ sky130_fd_sc_hd__dfstp_1
X_13764_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03263_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10976_ net672 _06469_ _06485_ net671 _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a221o_1
XFILLER_0_186_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09295__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15503_ clknet_leaf_42_wb_clk_i _01643_ _00311_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12715_ _06969_ _07238_ _06988_ _06949_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__or4b_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16483_ clknet_leaf_71_wb_clk_i net1550 _01291_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
X_13695_ net2137 _03217_ _03219_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__o21a_1
XANTENNA__11930__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15434_ clknet_leaf_37_wb_clk_i _01574_ _00242_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12646_ net266 net2001 net436 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ clknet_leaf_72_wb_clk_i _01505_ _00178_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[24\]
+ sky130_fd_sc_hd__dfstp_2
X_12577_ net252 net2045 net440 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14316_ net1209 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _05648_ _06116_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15296_ clknet_leaf_72_wb_clk_i _01440_ _00109_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold308 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold319 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14247_ net1173 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
X_11459_ net946 _06950_ _06954_ net604 vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__o211a_2
XFILLER_0_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_185_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09755__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ net1125 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XFILLER_0_194_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ _07375_ _07376_ _07415_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09507__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13303__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1019 team_02_WB.instance_to_wrap.ramload\[7\] vssd1 vssd1 vccd1 vccd1 net2381
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07621_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] _03337_ vssd1 vssd1 vccd1
+ vccd1 _03344_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_200_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ team_02_WB.instance_to_wrap.top.pc\[30\] vssd1 vssd1 vccd1 vccd1 _03293_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_191_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12001__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] net773 _04737_ _04738_
+ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a211o_1
XFILLER_0_173_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09038__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09153_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] net780 _04666_ _04667_
+ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03821_ _03822_ vssd1 vssd1
+ vccd1 vccd1 _03824_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_79_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11141__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A0 _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _04595_ _04597_ _04598_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__or4_1
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08035_ _03743_ _03751_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold820 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12671__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput80 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_1
Xinput91 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1131_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09746__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09210__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold886 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold897 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\] net825 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a22o_1
X_08937_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04293_ _04334_ vssd1
+ vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and3_2
XANTENNA__10108__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _04430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] _03532_ _03533_ vssd1 vssd1
+ vccd1 vccd1 _03542_ sky130_fd_sc_hd__and3_1
X_08799_ net1 net1038 vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nor2_1
X_10830_ net391 _06345_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__nor2_1
XANTENNA__10220__A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10761_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ _04334_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10292__A0 _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ net338 net2010 net557 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13480_ team_02_WB.START_ADDR_VAL_REG\[20\] _04260_ vssd1 vssd1 vccd1 vccd1 net204
+ sky130_fd_sc_hd__and2_1
X_10692_ _06201_ _06206_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__a21o_1
XANTENNA__09029__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ net325 net2110 net454 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13230__B1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10044__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15150_ net1158 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XANTENNA__09985__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ net313 net2240 net561 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__mux2_1
XANTENNA__11792__A0 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14101_ net1199 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11313_ net946 _06807_ _06814_ net604 vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__o211a_2
XANTENNA__12581__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15081_ net1253 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12293_ net308 net2255 net569 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
X_11244_ net409 _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__nor2_1
X_14032_ net1224 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XANTENNA__09737__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ _06180_ net653 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] net497
+ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] net927 net808 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15983_ clknet_leaf_43_wb_clk_i _02123_ _00791_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__B1 _06931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11925__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] net777 net773 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a22o_1
X_14934_ net1107 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
X_14865_ net1232 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
XANTENNA__13425__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13049__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ clknet_leaf_95_wb_clk_i _02723_ _01397_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_13816_ net1149 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
X_14796_ net1214 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XANTENNA__09268__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16535_ clknet_leaf_86_wb_clk_i _02662_ _01342_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_13747_ _03251_ net950 _03250_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959_ _06051_ _06060_ net394 vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11480__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16466_ clknet_leaf_70_wb_clk_i net1568 _01274_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
X_13678_ _03206_ _03209_ net1141 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_14_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15417_ clknet_leaf_123_wb_clk_i _01557_ _00225_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12629_ net1913 net327 net554 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16397_ clknet_leaf_99_wb_clk_i _02532_ _01205_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13221__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13275__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15415__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__C1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15348_ clknet_leaf_74_wb_clk_i _01488_ _00161_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09440__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12491__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 net140 vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ clknet_leaf_69_wb_clk_i _01423_ _00092_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 net121 vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net185 vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 _02616_ vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15565__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout607 _06281_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_4
X_09840_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] net895 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] net900 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\]
+ _05275_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a221o_1
XANTENNA__11835__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ _04262_ net1063 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10311__Y _05828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07604_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03325_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1 vccd1 _03327_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10040__A _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09259__A2 _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08584_ team_02_WB.instance_to_wrap.wb.curr_state\[2\] team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12666__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1081_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10274__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__A team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09205_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\] net797 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13212__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout604_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10026__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ _04630_ _04651_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__nand2_1
XANTENNA__09967__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\] net703 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08018_ _03696_ _03708_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__xnor2_2
Xhold650 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A _04284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold694 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] net738 _05484_ _05485_
+ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__a211o_1
XANTENNA__13279__B1 _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ _07492_ _07499_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__nand2_1
XANTENNA__09498__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11931_ net337 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\] net485 vssd1
+ vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10588__C _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14650_ net1096 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
X_11862_ net327 net2377 net492 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13601_ team_02_WB.instance_to_wrap.top.a1.row1\[10\] _03110_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[106\]
+ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10813_ _06319_ _06327_ net407 vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__mux2_1
XANTENNA__12576__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14581_ net1241 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
X_11793_ net321 net1925 net592 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ clknet_leaf_109_wb_clk_i _02460_ _01128_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15438__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10744_ team_02_WB.instance_to_wrap.top.pc\[14\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _06261_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16251_ clknet_leaf_32_wb_clk_i _02391_ _01059_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13203__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ team_02_WB.START_ADDR_VAL_REG\[3\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net217 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10675_ net789 _05669_ _06127_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o22a_4
X_15202_ net1247 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XFILLER_0_211_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12414_ net257 net2044 net454 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09958__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16182_ clknet_leaf_50_wb_clk_i _02322_ _00990_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13394_ net2615 net1013 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[23\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09422__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08630__A0 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ net1161 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
X_12345_ net238 net2310 net563 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_189_Left_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15064_ net1164 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
X_12276_ _04291_ net643 _07190_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or3_4
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14015_ net1115 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
X_11227_ net954 _06731_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_56_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11158_ _06544_ _06663_ net399 vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11508__X _07001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ _05580_ _05625_ net550 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__mux2_1
X_11089_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__inv_2
X_15966_ clknet_leaf_1_wb_clk_i _02106_ _00774_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09489__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917_ net1176 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_198_Left_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11296__A2 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ clknet_leaf_124_wb_clk_i _02037_ _00705_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14848_ net1106 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12486__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ net1089 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_193_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13171__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16518_ clknet_leaf_8_wb_clk_i _02652_ _01325_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10256__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09661__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16449_ clknet_leaf_44_wb_clk_i net1492 _01257_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07600__C team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09413__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15098__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08621__A0 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07609__A team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout404 _05900_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
Xfanout415 _05762_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_2
XANTENNA__08924__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 _07228_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08924__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09823_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\] net763 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\]
+ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a221o_1
Xfanout448 _07224_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_6
Xfanout459 _07220_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
XANTENNA__13346__A team_02_WB.instance_to_wrap.ramload\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09754_ net609 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__inv_2
X_08705_ _04308_ _04329_ net648 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__or3_2
X_09685_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] net803 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ _05189_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ team_02_WB.instance_to_wrap.top.a1.instruction\[2\] team_02_WB.instance_to_wrap.top.a1.instruction\[3\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[0\] team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_194_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout721_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _04180_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_202_Left_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout819_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13081__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\] net979 vssd1 vssd1 vccd1
+ vccd1 _04193_ sky130_fd_sc_hd__or2_1
XANTENNA__09652__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08860__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _05975_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09404__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09119_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] net866 vssd1 vssd1
+ vccd1 vccd1 _04636_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10391_ _05763_ net608 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_1__f_wb_clk_i_X clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12130_ net313 net2074 net468 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10970__A1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_211_Left_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ net299 net2596 net471 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XANTENNA__14640__A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold480 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ _06148_ _06234_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__xnor2_1
Xfanout960 _03261_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_2
X_15820_ clknet_leaf_126_wb_clk_i _01960_ _00628_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout971 net972 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 net985 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_2
XFILLER_0_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout993 _04427_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15751_ clknet_leaf_40_wb_clk_i _01891_ _00559_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12963_ team_02_WB.instance_to_wrap.top.pc\[8\] _05583_ vssd1 vssd1 vccd1 vccd1 _07483_
+ sky130_fd_sc_hd__nor2_1
Xhold1180 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14702_ net1083 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11914_ net267 net2387 net484 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__mux2_1
X_15682_ clknet_leaf_117_wb_clk_i _01822_ _00490_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12894_ _07380_ _07413_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09891__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14633_ net1214 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11845_ net258 net2123 net490 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10238__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14564_ net1134 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ net249 net1864 net594 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09643__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16303_ clknet_leaf_42_wb_clk_i _02443_ _01111_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13515_ _03072_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__nor2_1
X_10727_ _06168_ _06243_ _06167_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a21o_2
XANTENNA__08851__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14495_ net1115 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16234_ clknet_leaf_39_wb_clk_i _02374_ _01042_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13446_ _03036_ _03048_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__o21a_1
X_10658_ team_02_WB.instance_to_wrap.top.pc\[23\] _04494_ vssd1 vssd1 vccd1 vccd1
+ _06175_ sky130_fd_sc_hd__or2_1
Xclkload14 clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload25 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_6
XANTENNA__11570__A2_N net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload36 clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__11202__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16165_ clknet_leaf_30_wb_clk_i _02305_ _00973_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload47 clknet_leaf_92_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__inv_8
X_13377_ net2411 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[6\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10589_ net546 net391 net405 vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__or3_1
Xclkload58 clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__clkinv_8
Xclkload69 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__bufinv_16
X_15116_ net1105 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_12328_ net304 net2531 net565 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16096_ clknet_leaf_18_wb_clk_i _02236_ _00904_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15047_ net1230 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
X_12259_ net301 net1927 net573 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08906__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10713__A1 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_207_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15949_ clknet_leaf_48_wb_clk_i _02089_ _00757_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09470_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] net906 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09882__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08421_ _04117_ _04126_ _04123_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08352_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04059_ _04061_ _04062_ vssd1
+ vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09095__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08842__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ _03952_ _03994_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload8 clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11701__X _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1044_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10952__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1211_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout234 _07326_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
Xfanout245 net247 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 _03703_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_2
XANTENNA_fanout769_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] net913 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a22o_1
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10180__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07998_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03703_ vssd1 vssd1 vccd1
+ vccd1 _03721_ sky130_fd_sc_hd__xnor2_2
Xfanout289 net291 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
X_09737_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\] net787 net782 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09668_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] net767 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ _05169_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09873__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ net76 net1524 net957 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\] net812 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a22o_1
X_11630_ _05995_ _05996_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09086__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09625__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08833__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ net2298 net342 net638 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ team_02_WB.instance_to_wrap.ramaddr\[10\] net984 net966 _02999_ vssd1 vssd1
+ vccd1 vccd1 _01429_ sky130_fd_sc_hd__a22o_1
X_10512_ _04783_ _06028_ net536 _04776_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__o2bb2a_1
Xwire635 _04607_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14280_ net1111 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
X_11492_ net416 net666 _06569_ _06583_ _06983_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_21_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ net1417 _00012_ net939 _05855_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a22o_1
XANTENNA__13185__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ _04611_ _05959_ _04609_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__o21ba_1
XANTENNA_input65_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ _07484_ _07504_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__xor2_1
X_10374_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\] net918 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\]
+ _05886_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a221o_1
XANTENNA__10943__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15239__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12113_ net236 net2523 net466 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14370__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _07424_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__xor2_1
X_12044_ net242 net2237 net471 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11499__A2 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 _04327_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
X_15803_ clknet_leaf_30_wb_clk_i _01943_ _00611_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16783_ net1327 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_189_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13995_ net1124 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XFILLER_0_204_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11933__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15734_ clknet_leaf_21_wb_clk_i _01874_ _00542_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ team_02_WB.instance_to_wrap.top.pc\[17\] _06192_ vssd1 vssd1 vccd1 vccd1
+ _07466_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15665_ clknet_leaf_128_wb_clk_i _01805_ _00473_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12877_ _07388_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14616_ net1196 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
XANTENNA__09077__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ net327 net2361 net590 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_190_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15596_ clknet_leaf_126_wb_clk_i _01736_ _00404_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09616__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14547_ net1079 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_117_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11759_ net317 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\] net596 vssd1
+ vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08824__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14478_ net1076 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XANTENNA__10792__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload103 clknet_leaf_71_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__inv_8
Xclkload114 clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ clknet_leaf_125_wb_clk_i _02357_ _01025_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13429_ net1066 _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__nand2_2
X_16148_ clknet_leaf_3_wb_clk_i _02288_ _00956_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_188_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16079_ clknet_leaf_48_wb_clk_i _02219_ _00887_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08970_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] net739 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__a221o_1
X_07921_ _03605_ _03638_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_126_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07852_ _03304_ net329 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12004__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
X_07783_ _03303_ _03496_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11843__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09522_ _05016_ _05037_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10600__X _06117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08718__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09855__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _04962_ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nor2_8
XANTENNA_fanout252_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ _04111_ _04107_ _04099_ _04092_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__o2bb2a_1
X_09384_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\] net831 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a22o_1
XANTENNA__09068__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08335_ _04020_ _04038_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07618__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12674__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1259_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ _03958_ _03960_ _03938_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08197_ _03910_ _03912_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11178__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__A2 _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__X _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout886_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_144_Left_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1007 net1008 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\] net708 net701 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1018 team_02_WB.instance_to_wrap.top.ru.next_iready vssd1 vssd1 vccd1 vccd1
+ net1018 sky130_fd_sc_hd__clkbuf_2
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15799__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__B2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11753__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _04355_ _07123_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13780_ net1617 _03271_ _03273_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__a21oi_1
X_10992_ _06502_ _06503_ net412 vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__mux2_1
XANTENNA__11102__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09846__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ _06501_ _07254_ _06704_ _06730_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_153_Left_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15450_ clknet_leaf_53_wb_clk_i _01590_ _00258_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09059__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12662_ net325 net1950 net435 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ net1256 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_172_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _05831_ net657 _06113_ _05829_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_172_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12584__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ clknet_leaf_81_wb_clk_i _01521_ _00189_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08806__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16424__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ net312 net2363 net439 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__mux2_1
X_14332_ net1201 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11544_ net389 _07033_ _07034_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09178__B _04694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ net1208 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11475_ net670 _06957_ _06969_ net672 _06968_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__a221o_1
XANTENNA__11169__A1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16002_ clknet_leaf_119_wb_clk_i _02142_ _00810_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13214_ net629 net938 net1019 net1508 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a2bb2o_1
Xwire498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_8
X_10426_ _05167_ _05942_ _05168_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Left_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09231__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194_ net1183 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XANTENNA__11928__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _02908_ _02911_ net1027 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_150_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10357_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\] net785 net741 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a22o_1
X_13076_ _07363_ _07364_ _07428_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__and3_1
X_10288_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] net800 _05802_ _05803_
+ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a2111o_1
X_12027_ net298 net2501 net476 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10144__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16766_ net1310 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_171_Left_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13978_ net1095 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XANTENNA__09837__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15717_ clknet_leaf_28_wb_clk_i _01857_ _00525_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12929_ team_02_WB.instance_to_wrap.top.pc\[28\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _07449_ sky130_fd_sc_hd__nor2_1
X_16697_ net138 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15648_ clknet_leaf_17_wb_clk_i _01788_ _00456_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15579_ clknet_leaf_29_wb_clk_i _01719_ _00387_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ _03838_ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__and2_1
XANTENNA__09369__A _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08704__C _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ _03744_ _03750_ _03718_ _03732_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_180_Left_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09773__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10383__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__A team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _04462_ _04463_ _04467_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_168_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07904_ _03571_ _03600_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08884_ net11 net1032 net988 net2554 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10135__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07835_ _03546_ _03550_ _03557_ _03523_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a211o_1
XANTENNA__12669__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10978__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07766_ _03465_ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__and2_1
XANTENNA__09289__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] net898 net889 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07697_ _03403_ _03409_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a21o_1
XANTENNA__10843__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\] net717 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09367_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\] net715 _04880_ _04882_
+ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout801_A _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12596__A0 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08318_ _04000_ _04002_ _04018_ _04006_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09461__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\] net915 _04804_ _04805_
+ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a211o_1
XFILLER_0_191_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08249_ _03910_ _03925_ _03953_ _03960_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and4b_1
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14913__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _06188_ net653 _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a21o_1
XANTENNA__09213__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\] net764 _05717_ _05720_
+ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09285__Y _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ net374 _06437_ _06441_ net378 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10374__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10142_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] net703 _05655_ _05656_
+ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13248__B _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ net1213 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XANTENNA__13312__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10073_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\] net902 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a22o_1
XANTENNA__10126__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ net1254 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14881_ net1260 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12579__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__X _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16620_ clknet_leaf_90_wb_clk_i _02739_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13832_ net1155 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16551_ clknet_leaf_89_wb_clk_i _02675_ _01358_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_13763_ _03064_ net960 _03262_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__and3_1
X_10975_ net667 _06477_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15502_ clknet_leaf_47_wb_clk_i _01642_ _00310_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12714_ _07025_ _07237_ _07057_ _06996_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_48_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16482_ clknet_leaf_71_wb_clk_i net1490 _01290_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] _03217_ net1139 vssd1 vssd1
+ vccd1 vccd1 _03219_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15433_ clknet_leaf_111_wb_clk_i _01573_ _00241_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12645_ net258 net2288 net434 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ clknet_leaf_72_wb_clk_i _01504_ _00177_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_12576_ net238 net1935 net439 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315_ net1124 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
X_11527_ net419 _06636_ _06849_ net376 _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__a221o_2
XFILLER_0_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15295_ clknet_leaf_83_wb_clk_i _01439_ _00108_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13536__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ net1204 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
Xhold309 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ team_02_WB.instance_to_wrap.top.pc\[10\] net975 _06837_ _06953_ vssd1 vssd1
+ vccd1 vccd1 _06954_ sky130_fd_sc_hd__a211o_1
XANTENNA__09204__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10409_ _05513_ _05925_ _05514_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__o21a_1
X_14177_ net1258 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11389_ net998 _06887_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nor2_1
XANTENNA__10365__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ _07475_ _07512_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__xor2_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13303__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09923__Y _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ _07454_ _07530_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1009 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10798__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12489__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11393__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _03339_ _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_163_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1
+ _03292_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16749_ net1293 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09221_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\] net761 net721 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\] net715 _04668_ vssd1
+ vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09443__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08103_ _03821_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11141__B _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A1 _05510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] net925 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08034_ _03744_ _03750_ _03733_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_71_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput70 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
Xhold810 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xinput81 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_1
XFILLER_0_141_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold821 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
Xhold832 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold843 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 team_02_WB.instance_to_wrap.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net2249
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] net821 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\]
+ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout584_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04334_ vssd1 vssd1
+ vccd1 vccd1 _04453_ sky130_fd_sc_hd__nand2_1
XANTENNA__10108__A2 _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12399__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _04429_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout751_A _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _03532_ _03533_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1
+ vccd1 vccd1 _03541_ sky130_fd_sc_hd__a21oi_2
X_08798_ net2576 _04426_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07749_ _03432_ _03468_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__xor2_1
XANTENNA__10220__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13812__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ _04334_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09682__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09419_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\] net871 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a22o_1
XANTENNA__10292__A1 _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ _06198_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12430_ net322 net1835 net454 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13230__B2 _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12361_ net304 net2138 net562 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ net1239 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
X_11312_ _06192_ net652 _06809_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_134_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15080_ net1254 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12292_ net300 net2026 net570 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14031_ net1224 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
X_11243_ _06630_ _06746_ net398 vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10347__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__B1 _07001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _06227_ _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15247__Q team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\] net829 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\]
+ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a221o_1
XANTENNA__08960__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15982_ clknet_leaf_45_wb_clk_i _02122_ _00790_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14933_ net1225 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
X_10056_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\] net725 net721 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a22o_1
XANTENNA__12102__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14864_ net1256 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
XANTENNA__10411__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16603_ clknet_leaf_95_wb_clk_i _02722_ _01396_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13815_ net1138 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
X_14795_ net1124 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13746_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] _03019_ _03245_ vssd1
+ vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16534_ clknet_leaf_86_wb_clk_i _02661_ _01341_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_10958_ _06470_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09673__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13677_ _03198_ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or2_1
X_16465_ clknet_leaf_69_wb_clk_i net1447 _01273_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
X_10889_ _05809_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12628_ net2609 net321 net552 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__mux2_1
X_15416_ clknet_leaf_123_wb_clk_i _01556_ _00224_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09425__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16396_ clknet_leaf_80_wb_clk_i _02531_ _01204_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08779__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15347_ clknet_leaf_75_wb_clk_i _01487_ _00160_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_12559_ net304 net2335 net444 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15278_ clknet_leaf_66_wb_clk_i _01422_ _00091_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold106 _02572_ vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 net155 vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold128 _02617_ vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 team_02_WB.instance_to_wrap.ramstore\[2\] vssd1 vssd1 vccd1 vccd1 net1501
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ net1257 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_78_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10292__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] net891 _05272_ _05286_
+ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__a211o_1
XANTENNA__13288__B2 _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ _04287_ _04337_ _04342_ _04323_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_198_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1190 net1202 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_2
XANTENNA__12012__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] net998 vssd1 vssd1 vccd1
+ vccd1 _04281_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03325_ vssd1 vssd1 vccd1
+ vccd1 _03326_ sky130_fd_sc_hd__or2_1
X_08583_ team_02_WB.instance_to_wrap.wb.curr_state\[2\] team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11851__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11704__X _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09664__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13460__A1 team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07630__A team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout332_A _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\] net924 net920 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09416__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09135_ _04496_ _04650_ _04497_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12682__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1241_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] net719 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\]
+ _04582_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ _03675_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nand2_1
Xhold640 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10329__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold651 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold684 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\] net784 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a22o_1
XANTENNA__13279__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ net1419 _04441_ _04433_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\] net902 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ net325 net2078 net483 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_X clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ net323 net1683 net490 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
X_13600_ team_02_WB.instance_to_wrap.top.a1.row1\[18\] _03111_ _03116_ team_02_WB.instance_to_wrap.top.a1.row1\[122\]
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a22o_1
XANTENNA__11761__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10812_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__inv_2
X_14580_ net1241 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
XFILLER_0_200_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09655__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net320 net1838 net592 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _03085_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10743_ team_02_WB.instance_to_wrap.top.pc\[13\] team_02_WB.instance_to_wrap.top.pc\[12\]
+ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__and3_1
X_16250_ clknet_leaf_52_wb_clk_i _02390_ _01058_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13462_ team_02_WB.START_ADDR_VAL_REG\[2\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net214 sky130_fd_sc_hd__a21o_1
XANTENNA__16165__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input95_A wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ net994 _05693_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__and2_1
XANTENNA__13203__B2 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15201_ net1250 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
X_12413_ net251 net1829 net456 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_209_Right_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16181_ clknet_leaf_22_wb_clk_i _02321_ _00989_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12592__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ net2632 net1013 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[22\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15132_ net1158 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
X_12344_ net246 net2536 net561 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15063_ net1168 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
X_12275_ net348 net1834 net572 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
X_14014_ net1188 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
X_11226_ _04470_ _06713_ _06730_ net669 _06729_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__o221a_2
XANTENNA__09186__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11936__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__Y _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07645__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _06663_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] _04330_ net648 team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11088_ _05212_ _05980_ _06017_ _06020_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__o31a_1
X_15965_ clknet_leaf_11_wb_clk_i _02105_ _00773_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10039_ _05537_ _05555_ net969 vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__mux2_1
X_14916_ net1091 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
XANTENNA__09894__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15896_ clknet_leaf_121_wb_clk_i _02036_ _00704_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_160_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14847_ net1108 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14548__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14778_ net1095 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09646__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09110__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16517_ clknet_leaf_127_wb_clk_i _02651_ _01324_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16536__Q team_02_WB.instance_to_wrap.top.a1.row1\[58\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13729_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ _03017_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__and3_1
XFILLER_0_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16448_ clknet_leaf_43_wb_clk_i net1423 _01256_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07600__D team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16379_ clknet_leaf_86_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[3\] _01187_
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12007__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_2
X_09822_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\] net715 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a22o_1
XANTENNA__11846__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _07226_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_8
Xfanout449 _07224_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
X_09753_ _05259_ _05264_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__nor3_2
X_08704_ _04329_ net650 _04309_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__and3b_2
XANTENNA__13130__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\] net884 _05188_ _05200_
+ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a211o_1
XANTENNA__09885__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ team_02_WB.instance_to_wrap.top.a1.instruction\[4\] team_02_WB.instance_to_wrap.top.a1.instruction\[5\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04262_ vssd1 vssd1 vccd1 vccd1
+ _04264_ sky130_fd_sc_hd__nand4b_4
XANTENNA__12677__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08566_ _02814_ _04228_ _04226_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16188__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09637__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09101__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08497_ net1048 _04185_ _04191_ _04192_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout714_A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08743__X _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09118_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] net816 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\]
+ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a221o_1
X_10390_ _05763_ net608 vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09049_ net546 _04565_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ net311 net1804 net473 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold470 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net1832 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold481 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ net382 _06104_ _06513_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__a31o_2
Xhold492 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11756__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 _03233_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_2
Xfanout961 _03261_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout972 _04495_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_2
Xfanout994 net996 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13121__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15750_ clknet_leaf_8_wb_clk_i _01890_ _00558_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12962_ team_02_WB.instance_to_wrap.top.pc\[8\] _05583_ vssd1 vssd1 vccd1 vccd1 _07482_
+ sky130_fd_sc_hd__and2_1
XANTENNA__15405__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10486__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net257 net2203 net482 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__mux2_1
Xhold1181 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
X_14701_ net1122 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
Xhold1192 team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1 vccd1 vccd1 net2554
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12587__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ clknet_leaf_103_wb_clk_i _01821_ _00489_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12893_ _07379_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ net1105 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
X_11844_ net248 net1910 net491 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14563_ net1134 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
X_11775_ net253 net2018 net594 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XANTENNA__15260__Q team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ clknet_leaf_44_wb_clk_i _02442_ _01110_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_175_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10726_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] _04283_ _06169_ vssd1
+ vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__o21ai_1
X_13514_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__or4b_2
XFILLER_0_83_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ net1127 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13188__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13445_ _03033_ _02766_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__or3_1
X_16233_ clknet_leaf_112_wb_clk_i _02373_ _01041_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13212__A2_N net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657_ team_02_WB.instance_to_wrap.top.pc\[23\] _04491_ _04493_ vssd1 vssd1 vccd1
+ vccd1 _06174_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload15 clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload26 clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_6
XFILLER_0_140_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09197__A _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16164_ clknet_leaf_35_wb_clk_i _02304_ _00972_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload37 clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_6
X_13376_ team_02_WB.instance_to_wrap.ramload\[5\] net1011 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[5\] sky130_fd_sc_hd__and2_1
XANTENNA__09800__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10588_ _04458_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_58_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload48 clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_6
XFILLER_0_51_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload59 clknet_leaf_83_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_6
X_15115_ net1079 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ net298 net2283 net565 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__mux2_1
X_16095_ clknet_leaf_60_wb_clk_i _02235_ _00903_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_39_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_192_Right_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15046_ net1235 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XANTENNA__09159__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ net294 net1765 net574 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11209_ _06091_ _06095_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or2_1
X_12189_ net288 net2414 net576 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15948_ clknet_leaf_126_wb_clk_i _02088_ _00756_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09867__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12497__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15879_ clknet_leaf_38_wb_clk_i _02019_ _00687_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14278__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08420_ _04117_ _04126_ _04123_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08351_ _04061_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ _03995_ _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload9 clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12813__X _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1037_A _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10952__A2 _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10165__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09805_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\] net815 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a221o_1
Xfanout257 net260 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 _06564_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_1
X_07997_ _03716_ _03717_ _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__o211ai_1
Xfanout279 _06686_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout664_A _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13103__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\] net723 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a22o_1
XANTENNA__08738__X _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09667_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] net740 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\]
+ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__a221o_1
XANTENNA__11665__B1 _05533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_A _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1194_X net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ net77 net1420 net957 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
XANTENNA__12200__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _05109_ _05110_ _05112_ _05114_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__or4_1
XFILLER_0_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08549_ _04202_ _04203_ net651 net792 net1672 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11560_ net947 _07046_ _07050_ net605 vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__o211a_2
X_10511_ _05970_ _06027_ _05971_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire625 _05418_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11645__A2_N net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _05559_ net663 _06113_ _05557_ _06984_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire647 _05645_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_2
X_13230_ net1501 net1022 _02954_ _05807_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a22o_1
X_10442_ _05956_ _05958_ _04653_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11196__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ _07407_ _07408_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a21oi_1
X_10373_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\] net902 net804 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\]
+ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__a221o_1
XANTENNA__14651__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__A2 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ net247 net2458 net467 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input58_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _07366_ _07367_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__nand2b_1
X_12043_ net643 _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__nand2_1
XANTENNA__11339__X _06840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__X _05760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout780 _04367_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_4
Xfanout791 _04326_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
X_15802_ clknet_leaf_53_wb_clk_i _01942_ _00610_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16782_ net1326 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_204_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09849__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13994_ net1176 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XANTENNA__09313__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15733_ clknet_leaf_31_wb_clk_i _01873_ _00541_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11656__B1 _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ team_02_WB.instance_to_wrap.top.pc\[18\] _06190_ vssd1 vssd1 vccd1 vccd1
+ _07465_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_177_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ clknet_leaf_23_wb_clk_i _01804_ _00472_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12876_ _05695_ net500 vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14615_ net1186 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11827_ net321 net2354 net588 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
X_15595_ clknet_leaf_15_wb_clk_i _01735_ _00403_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_190_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11758_ net315 net1854 net598 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
X_14546_ net1178 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ _06224_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11689_ _05996_ _07129_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__nand2_1
X_14477_ net1120 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload104 clknet_leaf_72_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_126_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16216_ clknet_leaf_123_wb_clk_i _02356_ _01024_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13428_ team_02_WB.instance_to_wrap.top.lcd.currentState\[4\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ net962 vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13359_ team_02_WB.instance_to_wrap.ramload\[21\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[21\] sky130_fd_sc_hd__and2_1
X_16147_ clknet_leaf_52_wb_clk_i _02287_ _00955_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_188_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16078_ clknet_leaf_46_wb_clk_i _02218_ _00886_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ _03602_ _03639_ _03641_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13333__B1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15029_ net1261 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XANTENNA__10147__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire632_A _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _03548_ _03573_ _03572_ _03550_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__11895__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ _03503_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__nand2_1
XANTENNA__09390__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ _05016_ _05036_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08718__B _04346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\] net705 _04963_ _04966_
+ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12020__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08403_ net1645 net1008 net981 _04111_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09383_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\] net827 _04887_ _04899_
+ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a211o_1
XANTENNA__12808__X _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _03993_ _04045_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08265_ _03306_ _03974_ _03977_ _03966_ _03971_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a311o_1
XFILLER_0_116_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout412_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13291__A1_N _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08196_ _03910_ _03912_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12690__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14471__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09565__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout781_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A _04538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1148_X net2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10138__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 _03315_ vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1019 _00012_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09543__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13815__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11638__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\] net875 vssd1 vssd1
+ vccd1 vccd1 _05236_ sky130_fd_sc_hd__and2_1
X_10991_ _06294_ _06303_ net393 vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12730_ _06555_ _07253_ _06742_ _06768_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_195_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ net323 net1703 net434 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08066__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14400_ net1103 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ _05832_ _05905_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ net306 net2616 net441 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ clknet_leaf_83_wb_clk_i _01520_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11810__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11543_ net390 _06997_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__nand2_1
X_14331_ net1075 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XANTENNA__11070__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ net1120 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ _05925_ _06956_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13213_ net630 net937 net1021 net1415 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__a2bb2o_1
X_16001_ clknet_leaf_102_wb_clk_i _02141_ _00809_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ _05207_ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__or2_1
Xwire499 _05828_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_2
X_14193_ net1231 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XANTENNA__10377__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ _06259_ _06932_ net234 _02910_ net978 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__o32a_1
XANTENNA__09782__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] net765 net709 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\]
+ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13315__B1 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13075_ _07526_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10129__A0 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\] net914 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a22o_1
XANTENNA__12105__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ net309 net2052 net475 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XANTENNA__09534__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11944__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15893__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16765_ net1309 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
X_13977_ net1095 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
X_15716_ clknet_leaf_34_wb_clk_i _01856_ _00524_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12928_ _07446_ _07447_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__nand2_1
XANTENNA__10301__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16696_ net138 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11671__A_N _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15647_ clknet_leaf_61_wb_clk_i _01787_ _00455_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_157_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ net518 _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15578_ clknet_leaf_52_wb_clk_i _01718_ _00386_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10604__A1 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14529_ net1260 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ _03744_ _03750_ _03732_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10080__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10368__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__C1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09773__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07784__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13306__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ _04462_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__and2b_1
XANTENNA__12015__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__B team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11868__A0 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ _03593_ _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_4_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08883_ net12 net1032 net988 net2362 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_205_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11854__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _03520_ _03537_ _03554_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08729__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__B _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ _03441_ _03486_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_108_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09504_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] net927 net805 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\]
+ _05018_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07696_ _03414_ _03416_ _03418_ _03413_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_13__f_wb_clk_i_X clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09435_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\] net709 net681 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12685__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\] net691 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08317_ _04020_ _04021_ _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09297_ _04809_ _04810_ _04812_ _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09994__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _03930_ _03959_ _03963_ _03940_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o22a_1
XANTENNA__10071__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__X _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08179_ _03862_ _03889_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor2_2
X_10210_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\] net728 _05721_ _05723_
+ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_104_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11190_ net423 _06694_ _06695_ _06358_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09764__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\] net843 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\]
+ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a221o_1
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XANTENNA__09516__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\] net824 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\]
+ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a221o_1
XANTENNA__11764__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ net1263 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
X_14880_ net1104 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ net1150 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16550_ clknet_leaf_89_wb_clk_i _02674_ _01357_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10974_ _04734_ _06116_ _06467_ net664 _06486_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o221a_1
X_13762_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ clknet_leaf_48_wb_clk_i _01641_ _00309_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08077__C _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12713_ net672 _07032_ _07079_ _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_48_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16481_ clknet_leaf_69_wb_clk_i net1511 _01289_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
X_13693_ _03217_ _03218_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15432_ clknet_leaf_11_wb_clk_i _01572_ _00240_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ net249 net1817 net435 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ net245 net2168 net440 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15363_ clknet_leaf_72_wb_clk_i _01503_ _00176_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input80_X net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14314_ net1176 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
X_11526_ net397 _06939_ _07017_ net383 vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_152_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15294_ clknet_leaf_84_wb_clk_i _01438_ _00107_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11939__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13121__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14245_ net1114 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
X_11457_ net1000 _06952_ _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1
+ vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16691__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11011__A1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ _05558_ _05924_ _05557_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14176_ net1106 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XANTENNA__09755__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11388_ _06260_ _06886_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__or2_1
XANTENNA__08963__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ _05836_ _05855_ net968 vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__mux2_1
X_13127_ team_02_WB.instance_to_wrap.top.pc\[14\] net1023 _02896_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01495_ sky130_fd_sc_hd__a22o_1
XANTENNA__09507__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ _07433_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_X clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12009_ net643 _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__nand2_4
XANTENNA_wire428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16071__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__Y _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13067__A2 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07550_ net2323 vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__inv_2
X_16748_ net1292 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15639__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ clknet_leaf_65_wb_clk_i _02796_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09220_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] net733 net713 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11262__X _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16707__1349 vssd1 vssd1 vccd1 vccd1 net1349 _16707__1349/LO sky130_fd_sc_hd__conb_1
XFILLER_0_91_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\] net772 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08102_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03815_ _03816_ vssd1 vssd1
+ vccd1 vccd1 _03822_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] net891 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a22o_1
XANTENNA__10053__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11849__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ _03744_ _03754_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput60 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold800 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold811 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
Xmax_cap530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_1
XANTENNA__11538__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold833 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07628__A team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09746__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold844 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold855 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\] net923 net911 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1117_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04334_ vssd1 vssd1
+ vccd1 vccd1 _04452_ sky130_fd_sc_hd__and2_2
XANTENNA__12540__Y _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A _07214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08866_ net1382 net1038 net1037 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a21o_1
X_07817_ _03505_ _03535_ _03538_ _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_165_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08797_ team_02_WB.instance_to_wrap.top.pc\[0\] _04425_ _04357_ vssd1 vssd1 vccd1
+ vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout744_A _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_X clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_196_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12266__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _03468_ _03469_ vssd1 vssd1
+ vccd1 vccd1 _03471_ sky130_fd_sc_hd__or3_1
XFILLER_0_196_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09131__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ _03367_ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout911_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09418_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\] net903 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\]
+ _04929_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10690_ team_02_WB.instance_to_wrap.top.pc\[14\] _06197_ vssd1 vssd1 vccd1 vccd1
+ _06207_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09349_ _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10044__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12360_ net296 net2043 net561 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__mux2_1
XANTENNA__09985__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11759__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] net494 _06812_ _04263_ net496
+ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout999_X net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12291_ net292 net2163 net569 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__mux2_1
X_14030_ net1083 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XANTENNA__09198__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ _06745_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__inv_2
XANTENNA__09737__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _06181_ _06182_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__nand2b_1
X_10124_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\] net917 _05632_ _05633_
+ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a211o_1
XANTENNA_input40_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15981_ clknet_leaf_48_wb_clk_i _02121_ _00789_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] net784 _05561_ _05564_
+ _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a2111o_1
X_14932_ net1241 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_180_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09370__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14863_ net1219 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XANTENNA__15263__Q team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16602_ clknet_leaf_93_wb_clk_i _02721_ _01395_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13814_ net1138 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ net1188 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
XANTENNA__09122__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16533_ clknet_leaf_82_wb_clk_i net1019 _01340_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ _03245_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1
+ _03250_ sky130_fd_sc_hd__a31o_1
X_10957_ net408 _06044_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10283__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ clknet_leaf_69_wb_clk_i net1440 _01272_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13676_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _03208_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10888_ net405 _06350_ _06400_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_155_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15415_ clknet_leaf_115_wb_clk_i _01555_ _00223_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12627_ net2582 net317 net552 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16395_ clknet_leaf_87_wb_clk_i _02530_ _01203_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10035__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09928__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15346_ clknet_leaf_74_wb_clk_i _01486_ _00159_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_12558_ net297 net1917 net444 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ net418 _06356_ _06607_ _07000_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_20_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_max_cap542_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15277_ clknet_leaf_70_wb_clk_i _01421_ _00090_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 team_02_WB.instance_to_wrap.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net1469
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ net292 net2517 net557 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold118 net119 vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09189__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 team_02_WB.instance_to_wrap.ramstore\[22\] vssd1 vssd1 vccd1 vccd1 net1491
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228_ net1191 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ net1222 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_165_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12496__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _04328_ _04341_ _04345_ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1180 net1182 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__buf_4
X_08651_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] net998 vssd1 vssd1 vccd1
+ vccd1 _04280_ sky130_fd_sc_hd__nor2_4
Xfanout1191 net1194 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_198_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] team_02_WB.instance_to_wrap.top.a1.dataIn\[20\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1 vccd1 _03325_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_105_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11433__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09203_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] net822 net814 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\]
+ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout325_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ net969 _04650_ _04497_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09065_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\] net787 net779 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08016_ _03647_ _03660_ _03673_ _03645_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_116_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold630 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold652 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 team_02_WB.instance_to_wrap.top.a1.row1\[12\] vssd1 vssd1 vccd1 vccd1 net2025
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_A _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] net766 net720 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13279__A2 team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13095__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08918_ _04173_ _04209_ _04220_ net1010 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a32o_1
XANTENNA__12203__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\] net808 _05402_ _05414_
+ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__a211o_1
XANTENNA__09352__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08849_ net145 net1042 net1034 net1412 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XANTENNA__08418__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13823__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ net319 net1709 net490 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07821__A team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _06322_ _06326_ net372 vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__mux2_1
X_11791_ net313 net2200 net593 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _03073_ _03082_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__nor2_1
X_10742_ team_02_WB.instance_to_wrap.top.pc\[11\] _06258_ vssd1 vssd1 vccd1 vccd1
+ _06259_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13461_ team_02_WB.START_ADDR_VAL_REG\[1\] net1070 net1003 vssd1 vssd1 vccd1 vccd1
+ net203 sky130_fd_sc_hd__a21o_1
X_10673_ _06128_ _06189_ net790 _05625_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__13203__A2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ net1247 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
X_12412_ net254 net1900 net456 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16180_ clknet_leaf_4_wb_clk_i _02320_ _00988_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09958__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13392_ team_02_WB.instance_to_wrap.ramload\[21\] net1011 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[21\] sky130_fd_sc_hd__and2_1
XANTENNA_input88_A wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15131_ net1158 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
X_12343_ net240 net2199 net561 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10246__X _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15062_ net1263 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
X_12274_ net350 net2541 net572 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XANTENNA__15258__Q team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ _05974_ _06599_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__xor2_1
X_14013_ net1203 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
XANTENNA__09754__Y _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09591__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ net391 _06662_ _06661_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_208_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13717__B _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ net426 vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__inv_2
X_16706__1348 vssd1 vssd1 vccd1 vccd1 net1348 _16706__1348/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_147_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ _05948_ _05983_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12113__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15964_ clknet_leaf_19_wb_clk_i _02104_ _00772_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08099__A team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _05540_ _05549_ _05552_ _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__or4_2
X_14915_ net1136 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15895_ clknet_leaf_115_wb_clk_i _02035_ _00703_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11952__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ net1190 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14777_ net1098 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
X_11989_ net286 net2192 net478 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16516_ clknet_leaf_5_wb_clk_i _02650_ _01323_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_193_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13728_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03017_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a21o_1
XANTENNA__10256__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16447_ clknet_leaf_71_wb_clk_i net1466 _01255_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
X_13659_ net1374 net850 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11205__A1 _04284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16378_ clknet_leaf_86_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] _01186_
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15329_ clknet_leaf_42_wb_clk_i _01472_ _00142_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout406 _05900_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
Xfanout417 _05716_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_2
XANTENNA__09582__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\] net771 net746 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a22o_1
Xfanout439 _07226_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12023__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\] net715 _05266_ _05267_
+ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09334__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ _04283_ net789 vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__nand2_1
X_09683_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] net823 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout275_A _06740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ net1063 team_02_WB.instance_to_wrap.top.a1.instruction\[5\] team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__and4b_2
XANTENNA__07641__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__Y _06931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13362__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ team_02_WB.instance_to_wrap.top.a1.row1\[63\] _04225_ _04233_ _04183_ vssd1
+ vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout442_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08496_ team_02_WB.instance_to_wrap.top.a1.row1\[18\] net849 vssd1 vssd1 vccd1 vccd1
+ _04192_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12693__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09839__Y _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08860__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09117_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\] net922 net910 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1237_X net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ net972 _04564_ net544 vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold460 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11010_ net672 _06500_ _06501_ net671 _06521_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__a221o_1
Xhold482 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07816__A team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 _04532_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_8
Xfanout951 _03233_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_1
Xfanout962 _03027_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
Xfanout973 _04284_ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ team_02_WB.instance_to_wrap.top.pc\[10\] _05491_ vssd1 vssd1 vccd1 vccd1
+ _07481_ sky130_fd_sc_hd__and2_1
Xhold1160 team_02_WB.instance_to_wrap.top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 net2522
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11772__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1171 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ net1214 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1182 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net250 net2173 net484 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15680_ clknet_leaf_17_wb_clk_i _01820_ _00488_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1193 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08647__A team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _07383_ _07411_ _07381_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o21a_1
XANTENNA__07551__A team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ net1182 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
X_11843_ net252 net1991 net492 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11073__A _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10238__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14562_ net1130 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
XFILLER_0_200_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11774_ net239 net1799 net592 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
X_16301_ clknet_leaf_40_wb_clk_i _02441_ _01109_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _03072_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__nor2_1
X_10725_ _03293_ _06130_ _06241_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__o21ai_1
X_14493_ net1185 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XANTENNA__08851__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09478__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16232_ clknet_leaf_16_wb_clk_i _02372_ _01040_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13444_ _03028_ _03030_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10656_ team_02_WB.instance_to_wrap.top.pc\[24\] _06171_ vssd1 vssd1 vccd1 vccd1
+ _06173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_8
X_16163_ clknet_leaf_27_wb_clk_i _02303_ _00971_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10587_ _04458_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__and3_4
X_13375_ net2352 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[4\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12108__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload27 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__bufinv_16
Xclkload38 clknet_leaf_98_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_8
Xclkload49 clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_58_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15114_ net1102 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12326_ net310 net2141 net566 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__mux2_1
X_16094_ clknet_leaf_4_wb_clk_i _02234_ _00902_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11947__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__X _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ net1262 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
X_12257_ net287 net2539 net572 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11208_ _05944_ _05974_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__xnor2_1
X_12188_ net277 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\] net576 vssd1
+ vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11139_ _04951_ _06601_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__xnor2_1
X_15947_ clknet_leaf_14_wb_clk_i _02087_ _00755_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15878_ clknet_leaf_7_wb_clk_i _02018_ _00686_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09005__X _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14829_ net1121 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire508_A _05578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ _04047_ _04058_ _04049_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10229__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09095__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08281_ _03975_ _03994_ _03952_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08842__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13179__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12018__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13197__X _02953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16005__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09555__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net239 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
X_09804_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\] net831 net885 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__a22o_1
Xfanout247 _06372_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
Xfanout258 net260 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 _06626_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13639__C1 _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07996_ _03716_ _03717_ _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__o211a_1
XANTENNA__09307__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ net610 _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__nand2_1
XANTENNA__12688__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10997__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\] net755 net744 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ net78 team_02_WB.START_ADDR_VAL_REG\[15\] net956 vssd1 vssd1 vccd1 vccd1
+ _02643_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout824_A _04512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\] net833 net863 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_X net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _04199_ _04200_ net651 net792 net1455 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09086__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__X _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12276__X _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ net1064 _04176_ _03317_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__or3b_1
XANTENNA__08833__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10510_ _04866_ _06026_ _04862_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a21o_1
X_16705__1347 vssd1 vssd1 vccd1 vccd1 net1347 _16705__1347/LO sky130_fd_sc_hd__conb_1
XFILLER_0_147_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11490_ _05558_ net657 vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire626 _05332_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08654__D_N team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10441_ _04693_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__or2_1
XANTENNA__14932__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] net910 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13160_ net976 _07409_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11767__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12111_ net240 net2317 net468 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13091_ team_02_WB.instance_to_wrap.top.pc\[20\] net1025 _02866_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01501_ sky130_fd_sc_hd__a22o_1
XANTENNA__09546__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _06280_ _07201_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__nor2_2
Xhold290 team_02_WB.instance_to_wrap.top.a1.row2\[11\] vssd1 vssd1 vccd1 vccd1 net1652
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15801_ clknet_leaf_125_wb_clk_i _01941_ _00609_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout770 _04371_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout781 net784 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_8
X_16781_ net1325 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
Xfanout792 _04223_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_2
XFILLER_0_205_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13993_ net1216 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XANTENNA__11105__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12598__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15732_ clknet_leaf_14_wb_clk_i _01872_ _00540_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12944_ team_02_WB.instance_to_wrap.top.pc\[18\] _06190_ vssd1 vssd1 vccd1 vccd1
+ _07464_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_177_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15663_ clknet_leaf_48_wb_clk_i _01803_ _00471_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15271__Q team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ _07389_ _07393_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14614_ net1107 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11826_ net317 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\] net588 vssd1
+ vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
X_15594_ clknet_leaf_37_wb_clk_i _01734_ _00402_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09077__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14545_ net1231 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
X_11757_ net306 net2286 net599 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__mux2_1
XANTENNA__08824__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10092__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ team_02_WB.instance_to_wrap.top.pc\[20\] _06184_ vssd1 vssd1 vccd1 vccd1
+ _06225_ sky130_fd_sc_hd__xnor2_1
X_14476_ net1215 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
X_11688_ _07156_ _07161_ _07169_ _07173_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_155_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12908__A1 _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16215_ clknet_leaf_120_wb_clk_i _02355_ _01023_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11250__B _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ _03036_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__inv_2
Xclkload105 clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__inv_16
X_10639_ _04270_ _04288_ _04323_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__and3_1
XFILLER_0_180_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap1065 _03310_ vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09785__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16146_ clknet_leaf_54_wb_clk_i _02286_ _00954_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13358_ net2158 net1016 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[20\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_188_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12309_ _04291_ _04333_ _04452_ _06280_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__or4_2
X_16077_ clknet_leaf_50_wb_clk_i _02217_ _00885_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13289_ team_02_WB.instance_to_wrap.top.pc\[15\] net1054 _06830_ net933 vssd1 vssd1
+ vccd1 vccd1 _02994_ sky130_fd_sc_hd__a22o_1
X_15028_ net1230 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07850_ _03549_ net329 _03546_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire625_A _05418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07781_ _03303_ _03470_ net366 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__nand3_1
XANTENNA__13097__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__dlymetal6s2s_1
X_09520_ net970 net631 net543 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12301__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09451_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\] net721 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__a221o_1
X_08402_ _04102_ _04104_ _04108_ _04110_ _04097_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__a32o_2
X_09382_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] net929 net818 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\]
+ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a221o_1
XANTENNA__09068__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _03993_ _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10083__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ _03972_ _03979_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08195_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09528__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XANTENNA_fanout774_A _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08749__X _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _03677_ _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout941_A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\] net813 net905 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\]
+ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__a221o_1
XANTENNA__11638__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15695__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ net401 _06288_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09649_ net969 _05164_ _04497_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ net319 net1944 net434 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__mux2_1
XANTENNA_input105_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09059__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11611_ net379 _06502_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13260__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08806__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ net299 net1874 net440 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_67_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ net1087 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XANTENNA__10074__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11542_ _06046_ _06048_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_208_Left_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11070__B _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ net1224 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
X_11473_ _06966_ _06967_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16000_ clknet_leaf_18_wb_clk_i _02140_ _00808_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input70_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net632 net938 net1019 net1618 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a2bb2o_1
X_10424_ _05212_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and2_1
X_14192_ net1234 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XANTENNA__09231__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13143_ _07412_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__xnor2_1
X_10355_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\] net729 net681 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11069__Y _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13315__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\] net918 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__a22o_1
X_13074_ _07458_ _07459_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nor2_1
XANTENNA__10129__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__B1 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15266__Q team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12025_ net301 net1733 net476 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_183_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__X _06595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__A1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ net1308 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XANTENNA__12121__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ net1080 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XFILLER_0_205_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09298__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ clknet_leaf_9_wb_clk_i _01855_ _00523_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12927_ team_02_WB.instance_to_wrap.top.pc\[29\] _06140_ vssd1 vssd1 vccd1 vccd1
+ _07447_ sky130_fd_sc_hd__or2_1
X_16695_ net138 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11960__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15646_ clknet_leaf_5_wb_clk_i _01786_ _00454_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12858_ net789 _04417_ _06127_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_85_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ net252 net1823 net589 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15577_ clknet_leaf_121_wb_clk_i _01717_ _00385_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12789_ _06344_ _06398_ _06446_ _06477_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__and4_1
XFILLER_0_145_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10065__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528_ net1081 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11262__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14459_ net1087 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09758__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08570__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12804__B _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ clknet_leaf_100_wb_clk_i _02269_ _00937_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08951_ _04463_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__nor2_1
XANTENNA__07617__C team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07902_ _03554_ _03570_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08882_ net14 net1030 net987 net2158 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__o22a_1
XFILLER_0_209_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_205_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09930__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07833_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__inv_2
X_16704__1346 vssd1 vssd1 vccd1 vccd1 net1346 _16704__1346/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12031__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _03461_ _03462_ _03437_ _03441_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09289__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09503_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\] net799 net863 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a221o_1
XANTENNA__13319__A1_N _07183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ _03380_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__and2b_1
XANTENNA__11870__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1097_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _04948_ _04949_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__nand2b_2
XANTENNA__10843__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09365_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] net775 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\]
+ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XANTENNA__10339__X _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1264_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10056__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ _04028_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\] net920 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ _04803_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a221o_1
XANTENNA__09461__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08247_ _03938_ _03958_ _03960_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _03321_ _03896_ net2125 net1007 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09213__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12206__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10140_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] net778 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a22o_1
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
X_10071_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\] net918 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a22o_1
X_13830_ net1150 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13761_ net2584 net960 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__and2b_1
XFILLER_0_168_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _04778_ net662 _06484_ net795 vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_168_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11780__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14657__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15500_ clknet_leaf_2_wb_clk_i _01640_ _00308_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12712_ _07100_ _07113_ _07129_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__and3_1
XANTENNA__10295__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16480_ clknet_leaf_71_wb_clk_i net1481 _01288_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
X_13692_ net1603 _03216_ net1066 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_48_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15431_ clknet_leaf_38_wb_clk_i _01571_ _00239_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12643_ net252 net2244 net436 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ clknet_leaf_82_wb_clk_i _01502_ _00175_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_12574_ net242 net2592 net440 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08942__X _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09452__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14313_ net1221 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11525_ net407 _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_152_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15293_ clknet_leaf_83_wb_clk_i _01437_ _00106_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13536__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ net1093 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
X_11456_ _06258_ _06951_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09204__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ _05918_ _05923_ _05604_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11011__A2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12116__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14175_ net1108 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
X_11387_ team_02_WB.instance_to_wrap.top.pc\[12\] _06259_ team_02_WB.instance_to_wrap.top.pc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_185_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ net976 _07417_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__o31ai_1
X_10338_ _05845_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__or2_4
XANTENNA__10770__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11955__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ net535 _06150_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__xnor2_1
X_10269_ _05740_ _05785_ net550 vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__mux2_1
XANTENNA__09912__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _07190_ _07201_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_163_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_187_Right_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16747_ team_02_WB.instance_to_wrap.top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 net178
+ sky130_fd_sc_hd__clkbuf_1
X_13959_ net1169 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_93_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10286__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16678_ clknet_leaf_65_wb_clk_i _02795_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15240__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13224__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15629_ clknet_leaf_48_wb_clk_i _01769_ _00437_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09150_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\] net754 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a22o_1
XANTENNA__09979__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ _03815_ _03816_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1
+ vccd1 vccd1 _03821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09081_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\] net830 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ _04590_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08032_ _03711_ _03753_ _03706_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__a21o_1
Xinput50 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
Xhold801 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold812 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
Xhold823 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap542 _04672_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_4
Xhold834 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xinput94 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_1
XANTENNA__12026__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold845 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] net817 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__a221o_1
XANTENNA__11865__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ team_02_WB.instance_to_wrap.top.a1.row1\[101\] _03319_ vssd1 vssd1 vccd1
+ vccd1 _02515_ sky130_fd_sc_hd__or2_1
XANTENNA__10622__X _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1012_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13365__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ net138 _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout472_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] _03470_ _03506_ vssd1 vssd1
+ vccd1 vccd1 _03539_ sky130_fd_sc_hd__or3_1
X_08796_ _04423_ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12696__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ _03468_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout737_A _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10277__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07678_ _03393_ _03394_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _03364_ vssd1
+ vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09682__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11172__Y _06679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09417_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\] net830 net925 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\]
+ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13215__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10029__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ _04863_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08762__X _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09279_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\] net703 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\]
+ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a221o_1
X_11310_ _06811_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__inv_2
XANTENNA__07819__A team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12290_ net286 net2395 net569 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11529__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _06688_ _06744_ net370 vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__mux2_1
XANTENNA__10201__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _06677_ _06678_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _05635_ _05636_ _05638_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15980_ clknet_leaf_126_wb_clk_i _02120_ _00788_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ net1086 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
X_10054_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\] net701 _05565_ _05567_
+ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_180_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10504__A1 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ net1083 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XANTENNA__08937__X _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16601_ clknet_leaf_93_wb_clk_i _02720_ _01394_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13813_ net1155 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
X_14793_ net1210 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07560__Y _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16532_ clknet_leaf_80_wb_clk_i _00007_ _01339_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13744_ net2167 _03247_ _03249_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__o21a_1
X_10956_ _06467_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09673__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16463_ clknet_leaf_69_wb_clk_i net1458 _01271_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13675_ _03206_ _03207_ net1139 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10887_ net382 _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ clknet_leaf_21_wb_clk_i _01554_ _00222_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ net1982 net312 net554 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_159_Left_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16394_ clknet_leaf_80_wb_clk_i _02529_ _01202_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09425__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15345_ clknet_leaf_73_wb_clk_i _01485_ _00158_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_12557_ net308 net2446 net442 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XANTENNA__11232__A2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16703__1345 vssd1 vssd1 vccd1 vccd1 net1345 _16703__1345/LO sky130_fd_sc_hd__conb_1
X_11508_ net418 _06607_ _06608_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__a31o_1
X_15276_ clknet_leaf_84_wb_clk_i _01420_ _00089_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12488_ net284 net2534 net556 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
Xhold108 team_02_WB.instance_to_wrap.ramstore\[7\] vssd1 vssd1 vccd1 vccd1 net1470
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14227_ net1072 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
Xhold119 _02615_ vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ net948 _06931_ _06935_ net607 vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__o211a_2
XFILLER_0_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14158_ net1076 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13109_ team_02_WB.instance_to_wrap.top.pc\[17\] net1023 _02881_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01498_ sky130_fd_sc_hd__a22o_1
XANTENNA__11538__X _07030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ net1216 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_168_Left_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15606__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1170 net1171 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_4
X_08650_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net1060 net997 _04277_
+ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__and4_1
Xfanout1192 net1194 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_198_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07601_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_105_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ team_02_WB.instance_to_wrap.wb.curr_state\[0\] _04242_ vssd1 vssd1 vccd1
+ vccd1 _04243_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09664__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\] net830 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09416__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _04640_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__or2_4
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout318_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09064_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] net767 _04571_ _04573_
+ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10982__A1 _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08015_ _03736_ _03734_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10982__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold620 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold653 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\] net757 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a22o_1
X_08917_ net1404 _04440_ net930 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
X_09897_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] net926 net922 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\]
+ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a221o_1
XANTENNA__13684__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ net1487 net1043 net1035 team_02_WB.instance_to_wrap.ramstore\[16\] vssd1
+ vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
X_08779_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\] net761 net745 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10810_ _06324_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11790_ net304 net2574 net595 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XANTENNA__09655__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ team_02_WB.instance_to_wrap.top.pc\[10\] team_02_WB.instance_to_wrap.top.pc\[9\]
+ _06257_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and3_1
XANTENNA__08863__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ team_02_WB.EN_VAL_REG net1069 net1003 _03060_ vssd1 vssd1 vccd1 vccd1 net192
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_36_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ net995 _05669_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09407__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08615__A0 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12411_ net237 net2066 net454 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ net2158 net1013 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[20\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08652__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15130_ net1158 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _04292_ net643 _07193_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10973__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15061_ net1253 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
X_12273_ net363 net2196 net572 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15629__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ net1192 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
X_11224_ net654 _06720_ _06728_ net794 _06725_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__o221a_1
XANTENNA__08918__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09040__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _04970_ net387 _06097_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_56_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13717__C net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net698 _05616_ _05621_
+ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a2111oi_4
XTAP_TAPCELL_ROW_147_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ net2100 net262 net639 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
X_15963_ clknet_leaf_29_wb_clk_i _02103_ _00771_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_147_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10037_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] net818 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\]
+ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a221o_1
X_14914_ net1153 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
X_15894_ clknet_leaf_49_wb_clk_i _02034_ _00702_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09894__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14845_ net1205 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15006__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14776_ net1198 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
X_11988_ net272 net2435 net479 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XANTENNA__09646__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16515_ clknet_leaf_127_wb_clk_i _02649_ _01322_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13727_ net950 _03237_ _03238_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__and3_1
X_10939_ net380 _06449_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__or2_1
XANTENNA__08854__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16446_ clknet_leaf_45_wb_clk_i net1416 _01254_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
X_13658_ net1371 _04134_ net850 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ net1814 net238 net555 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16377_ clknet_leaf_85_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[1\] _01185_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13589_ _03289_ team_02_WB.instance_to_wrap.top.lcd.nextState\[2\] _03142_ _03122_
+ team_02_WB.instance_to_wrap.top.a1.row2\[9\] vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15328_ clknet_leaf_72_wb_clk_i _01471_ _00141_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15259_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[18\]
+ _00072_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12166__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14580__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09031__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
X_09820_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] net775 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a22o_1
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_2
XANTENNA__12304__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\] net763 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a22o_1
X_08702_ net994 net791 vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__nor2_1
XANTENNA__10900__X _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\] net924 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09885__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ team_02_WB.instance_to_wrap.top.a1.instruction\[0\] team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 _04262_
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_87_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout268_A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09098__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _04227_ _04229_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_178_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09637__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08845__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08495_ team_02_WB.instance_to_wrap.top.a1.data\[10\] net958 _04190_ vssd1 vssd1
+ vccd1 vccd1 _04191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout435_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1177_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout602_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\] net824 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09047_ _04546_ _04558_ _04561_ _04563_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__nor4_2
Xhold450 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold483 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12214__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold494 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10183__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 _04433_ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 _04532_ vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_4
X_09949_ net514 _05464_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and2_1
Xfanout952 _04499_ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_2
Xfanout963 _03027_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_205_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net975 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
Xfanout985 _02956_ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 _04282_ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ team_02_WB.instance_to_wrap.top.pc\[10\] _05491_ vssd1 vssd1 vccd1 vccd1
+ _07480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1150 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09876__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702__1344 vssd1 vssd1 vccd1 vccd1 net1344 _16702__1344/LO sky130_fd_sc_hd__conb_1
Xhold1161 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ net252 net2425 net484 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__mux2_1
Xhold1172 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ _07384_ _07410_ _07385_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__o21ba_1
Xhold1194 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
X_14630_ net1213 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11842_ net236 net2289 net490 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14561_ net1259 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
XANTENNA__11073__B _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07639__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ net247 net1942 net594 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16300_ clknet_leaf_126_wb_clk_i _02440_ _01108_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13512_ team_02_WB.instance_to_wrap.top.pad.keyCode\[6\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_175_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _06132_ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_175_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ net1192 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
X_16231_ clknet_leaf_39_wb_clk_i _02371_ _01039_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13443_ _03033_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__nor2_1
X_10655_ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__inv_2
XFILLER_0_192_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11199__A1 _04469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16162_ clknet_leaf_118_wb_clk_i _02302_ _00970_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload17 clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_8
X_13374_ net2572 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[3\]
+ sky130_fd_sc_hd__and2_1
X_10586_ net667 _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nor2_1
XANTENNA__15269__Q team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload28 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_8
XANTENNA__09800__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload39 clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_58_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15113_ net1103 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
X_12325_ net300 net2547 net565 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__mux2_1
X_16093_ clknet_leaf_12_wb_clk_i _02233_ _00901_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15044_ net1260 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
X_12256_ net275 net2258 net573 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11207_ net1777 net289 net638 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12187_ net282 net2319 net578 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__mux2_1
XANTENNA__12124__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ net656 _06637_ _06642_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11963__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ net398 _06578_ _06575_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__a21oi_4
X_15946_ clknet_leaf_39_wb_clk_i _02086_ _00754_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09867__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ clknet_leaf_30_wb_clk_i _02017_ _00685_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14828_ net1209 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_176_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09619__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14759_ net1182 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08280_ _03952_ _03975_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__X _04538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13179__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ clknet_leaf_64_wb_clk_i net1502 _01237_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10608__A _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09252__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12034__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\] net909 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\]
+ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout237 net239 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11362__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 _06498_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
X_07995_ _03716_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nor2_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_1
XFILLER_0_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ net970 _05250_ net543 vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10997__B _06508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] net731 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\]
+ _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout552_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08616_ net79 net1532 _04261_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09596_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] net918 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.row1\[111\]
+ net793 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XANTENNA__08818__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout817_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08478_ _00017_ _03317_ _04175_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12209__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__A _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire627 _05289_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ _04630_ _04651_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08770__X _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\] net813 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ _05883_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12110_ net643 _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__nand2_1
X_13090_ _04280_ _02864_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11445__A1_N net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ net346 net2455 net474 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__mux2_1
Xhold280 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11783__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 _04374_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_144_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15800_ clknet_leaf_120_wb_clk_i _01940_ _00608_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout771 _04371_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_8
Xfanout782 net784 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_8
X_16780_ net1324 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
X_13992_ net1113 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
Xfanout793 _04223_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08658__A _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15731_ clknet_leaf_59_wb_clk_i _01871_ _00539_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12943_ team_02_WB.instance_to_wrap.top.pc\[19\] _06188_ vssd1 vssd1 vccd1 vccd1
+ _07463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ clknet_leaf_46_wb_clk_i _01802_ _00470_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12874_ _05742_ net608 vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_29_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14613_ net1257 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
X_11825_ net315 net1949 net590 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
X_15593_ clknet_leaf_116_wb_clk_i _01733_ _00401_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08809__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14544_ net1225 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ net299 net2439 net598 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
XANTENNA__09482__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ team_02_WB.instance_to_wrap.top.pc\[19\] _06186_ _06223_ vssd1 vssd1 vccd1
+ vccd1 _06224_ sky130_fd_sc_hd__a21oi_1
X_14475_ net1100 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
X_11687_ _04569_ _04589_ _04608_ _07170_ _07172_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__o311a_1
XFILLER_0_181_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12119__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16214_ clknet_leaf_49_wb_clk_i _02354_ _01022_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13426_ _03289_ net962 _03035_ net1145 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_155_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10638_ _04272_ _04277_ net1060 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13030__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload106 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_16
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16145_ clknet_leaf_128_wb_clk_i _02285_ _00953_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11958__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ team_02_WB.instance_to_wrap.ramload\[19\] net1016 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[19\] sky130_fd_sc_hd__and2_1
X_10569_ net407 _06078_ _06083_ net380 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12308_ net349 net1969 net568 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__mux2_1
Xmax_cap949 _03355_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__buf_1
XFILLER_0_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_188_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16076_ clknet_leaf_126_wb_clk_i _02216_ _00884_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13288_ net1482 net983 net965 _02993_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15027_ net1234 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12239_ net1664 net356 net614 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XANTENNA__10147__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_207_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07780_ _03303_ net366 _03470_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__a21o_1
XANTENNA_wire520_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_15929_ clknet_leaf_124_wb_clk_i _02069_ _00737_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\] net733 net685 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__a22o_1
X_08401_ _04096_ _04098_ _04094_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a21o_1
X_09381_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\] net885 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08332_ _03306_ _03990_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload72_A clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08263_ _03306_ _03974_ _03977_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12029__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09225__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ _03823_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11868__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16701__1343 vssd1 vssd1 vccd1 vccd1 net1343 _16701__1343/LO sky130_fd_sc_hd__conb_1
XFILLER_0_6_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13649__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13368__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10138__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11335__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12699__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16272__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13384__A team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10801__A _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ _03668_ _03699_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08478__A _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09717_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\] net917 net801 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11638__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16695__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _04496_ _05164_ _04497_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08765__X _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10310__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\] net753 _05094_ _05095_
+ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11610_ _05999_ _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12590_ net309 net2033 net439 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__mux2_1
XANTENNA__09464__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _05912_ _05916_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_122_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14260_ net1241 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XANTENNA__09216__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ net663 _06956_ _06965_ net655 _06958_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__o221a_1
X_13211_ _04990_ net936 net1020 net1422 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_137_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11778__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _05935_ _05938_ _05252_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__o21a_1
X_14191_ net1196 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10377__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ _07379_ _07380_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nand2_1
X_10354_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\] net781 net773 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\]
+ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a221o_1
XANTENNA_input63_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09519__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11079__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13315__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13073_ net1027 _02851_ net1025 team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1
+ vccd1 vccd1 _01504_ sky130_fd_sc_hd__a2bb2o_1
X_10285_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\] net808 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__a221o_1
X_12024_ net294 net1918 net476 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_131_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10270__X _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12402__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13079__A1 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_164_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13079__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16763_ net1307 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
X_13975_ net1169 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
X_15714_ clknet_leaf_116_wb_clk_i _01854_ _00522_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12926_ team_02_WB.instance_to_wrap.top.pc\[29\] _06140_ vssd1 vssd1 vccd1 vccd1
+ _07446_ sky130_fd_sc_hd__nand2_1
X_16694_ net138 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10301__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10857__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15645_ clknet_leaf_10_wb_clk_i _01785_ _00453_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12857_ _05355_ _06205_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ net236 net2327 net591 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_140_Left_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12788_ _06508_ _06541_ _06573_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__and3_1
XANTENNA__09455__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15576_ clknet_leaf_121_wb_clk_i _01716_ _00384_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10065__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09012__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14527_ net1108 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11739_ net243 net1957 net598 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09207__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14458_ net1087 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13409_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or4b_1
X_14389_ net1257 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16128_ clknet_leaf_110_wb_clk_i _02268_ _00936_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08950_ _04276_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__nand2_4
XANTENNA__13306__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16059_ clknet_leaf_32_wb_clk_i _02199_ _00867_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11317__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ _03562_ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_168_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ net15 net1032 net988 net2527 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ _03520_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12312__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10621__A team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07763_ _03461_ _03462_ _03437_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09502_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] net821 net817 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08497__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07694_ _03345_ _03347_ _03361_ _03351_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ _04928_ _04947_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout250_A _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout348_A _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09364_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\] net759 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09446__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08315_ _04000_ _04002_ _04018_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09295_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\] net903 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\]
+ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14763__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1257_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08246_ _03961_ _03959_ _03932_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13379__A team_02_WB.instance_to_wrap.ramload\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08177_ _03888_ _03893_ _03862_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15367__Q team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10764__C1 team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__clkbuf_4
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_11_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
X_10070_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\] net874 net863 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ _05586_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12222__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _03065_ _03258_ _03259_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o211a_1
X_10972_ _06029_ _06467_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09685__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12711_ _06125_ _07234_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__nor2_1
X_13691_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\] _03216_ vssd1 vssd1 vccd1
+ vccd1 _03217_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12642_ net236 net2415 net434 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__mux2_1
X_15430_ clknet_leaf_9_wb_clk_i _01570_ _00238_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09437__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ clknet_leaf_82_wb_clk_i _01501_ _00174_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_12573_ net642 _07207_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__nand2_8
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11524_ _06978_ _07015_ net367 vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__mux2_1
X_14312_ net1111 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
X_15292_ clknet_leaf_70_wb_clk_i _01436_ _00105_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08671__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14243_ net1134 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13536__A2 _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ team_02_WB.instance_to_wrap.top.pc\[9\] _06257_ team_02_WB.instance_to_wrap.top.pc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14174_ net1189 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ team_02_WB.instance_to_wrap.top.pc\[12\] _06205_ _06203_ vssd1 vssd1 vccd1
+ vccd1 _06885_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_185_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ net229 _02893_ _06861_ net232 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__o2bb2a_1
X_10337_ _05847_ _05849_ _05851_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08963__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ _06560_ net235 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__nor2_1
XANTENNA__08610__S _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10268_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] net648 _05784_ vssd1
+ vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a21o_1
X_12007_ net346 net2552 net478 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15009__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12132__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ net969 _05695_ _05714_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11971__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16746_ net1291 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_205_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09676__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16700__1342 vssd1 vssd1 vccd1 vccd1 net1342 _16700__1342/LO sky130_fd_sc_hd__conb_1
X_13958_ net1249 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_200_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09140__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12909_ _07364_ _07428_ _07363_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__a21oi_1
X_16677_ clknet_leaf_65_wb_clk_i _02794_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13889_ net1250 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XANTENNA__11272__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ clknet_leaf_124_wb_clk_i _01768_ _00436_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09013__Y _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13224__B2 _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ clknet_leaf_38_wb_clk_i _01699_ _00367_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ _03818_ _03819_ _03799_ _03817_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o2bb2a_1
X_09080_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\] net920 net912 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\]
+ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_204_Right_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ _03740_ _03741_ _03743_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__o31a_1
Xinput40 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13199__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12307__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap510 _05533_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold802 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xinput62 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_2
Xmax_cap521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_2
Xinput73 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput84 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
Xhold813 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_1
Xhold835 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold846 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold868 team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net2230
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\] net893 net889 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a22o_1
Xhold879 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12831__A _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__A team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net1437 _04451_ net930 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_A _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net1503 net1039 net1037 team_02_WB.instance_to_wrap.ramstore\[0\] vssd1 vssd1
+ vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
X_07815_ _03532_ _03533_ _03507_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08795_ net548 _04422_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nand2_1
XANTENNA__14758__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03461_ _03462_ vssd1 vssd1
+ vccd1 vccd1 _03469_ sky130_fd_sc_hd__and3_1
XANTENNA__09667__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09131__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _03364_ _03396_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__xor2_2
XFILLER_0_177_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08475__B team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09416_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] net900 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09419__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13215__B2 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ net533 _04861_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09858__Y _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\] net727 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ _03916_ _03926_ _03918_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10085__X _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12217__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _06333_ _06336_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__nand2_1
XANTENNA__09198__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ net837 _06658_ _06660_ net669 vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__o22a_1
XANTENNA__10960__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\] net919 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\]
+ _05634_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\] net785 _05568_ _05569_
+ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a211o_1
X_14930_ net1184 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_180_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15408__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1123 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XANTENNA__11791__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ clknet_leaf_90_wb_clk_i _02719_ _01393_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13812_ net1142 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
XANTENNA__09658__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14792_ net1111 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XANTENNA__09122__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16531_ clknet_leaf_84_wb_clk_i net1373 _01338_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10955_ _04777_ _05954_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__and2b_1
X_13743_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] _03247_ net951 vssd1
+ vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_211_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16462_ clknet_leaf_66_wb_clk_i net1430 _01270_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10886_ net407 _06400_ _06352_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08953__X _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15413_ clknet_leaf_32_wb_clk_i _01553_ _00221_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12625_ net2358 net305 net553 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16393_ clknet_leaf_99_wb_clk_i _02528_ _01201_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12556_ net303 net2271 net444 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15344_ clknet_leaf_73_wb_clk_i _01484_ _00157_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08605__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ _06087_ _06820_ _06999_ net383 vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a22o_1
X_12487_ net273 net2338 net559 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__mux2_1
XANTENNA__12127__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ clknet_leaf_84_wb_clk_i _01419_ _00088_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold109 _02569_ vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09189__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11438_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _06833_ _06934_ vssd1 vssd1
+ vccd1 vccd1 _06935_ sky130_fd_sc_hd__a21o_1
X_14226_ net1178 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11966__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ net1122 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
X_11369_ _06062_ _06064_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_210_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap528_A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ _02878_ _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__o21ai_1
X_14088_ net1112 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_165_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13039_ _07449_ _07450_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and2b_1
XANTENNA__09897__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__buf_4
XANTENNA__09361__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1171 net1265 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_8
Xfanout1182 net1187 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_198_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_2
X_07600_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] team_02_WB.instance_to_wrap.top.a1.dataIn\[26\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__or4_1
X_08580_ team_02_WB.instance_to_wrap.Wen team_02_WB.instance_to_wrap.Ren vssd1 vssd1
+ vccd1 vccd1 _04242_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_105_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09649__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16729_ net1357 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] net900 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_56_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09132_ _04642_ _04644_ _04646_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08624__A1 team_02_WB.START_ADDR_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10617__Y _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\] net744 _04574_ _04576_
+ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_44_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12037__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08014_ _03736_ _03734_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__and2b_1
XANTENNA__10982__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold610 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 team_02_WB.instance_to_wrap.ramaddr\[12\] vssd1 vssd1 vccd1 vccd1 net1983
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_116_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11876__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold654 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold665 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold676 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] net732 _05471_ _05474_
+ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout582_A _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ _04173_ _04206_ _04217_ net1009 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__a32o_1
XANTENNA__09888__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] net890 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1008_X net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net147 net1044 net1036 net1434 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ net847 _04363_ _04364_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__and3_1
XANTENNA__09104__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ _03416_ _03449_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ team_02_WB.instance_to_wrap.top.pc\[8\] _06256_ vssd1 vssd1 vccd1 vccd1 _06257_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08773__X _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ net789 _05580_ _06127_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12410_ net246 net2007 net457 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13390_ team_02_WB.instance_to_wrap.ramload\[19\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[19\] sky130_fd_sc_hd__and2_1
XANTENNA__09812__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12341_ net346 net2605 net564 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15060_ net1251 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
X_12272_ net354 net2190 net574 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14011_ net1082 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
XANTENNA__11786__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11639__X _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10186__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A2 _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07565__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net371 _06604_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__or2_1
XANTENNA__09591__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10105_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\] net712 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__a22o_1
X_15962_ clknet_leaf_18_wb_clk_i _02102_ _00770_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11085_ net606 _06589_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_147_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09879__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14913_ net1261 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
X_10036_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\] net925 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__a22o_1
X_15893_ clknet_leaf_40_wb_clk_i _02033_ _00701_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12410__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14844_ net1201 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08396__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14775_ net1186 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11987_ net290 net1782 net481 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ clknet_leaf_5_wb_clk_i _02648_ _01321_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13726_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03017_ vssd1 vssd1 vccd1
+ vccd1 _03238_ sky130_fd_sc_hd__nand2_1
X_10938_ net424 _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10110__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16445_ clknet_leaf_71_wb_clk_i net1509 _01253_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10869_ net389 _06050_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a21oi_1
X_13657_ net1390 _04143_ net850 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11550__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12608_ net1891 net246 net553 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16376_ clknet_leaf_86_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[0\] _01184_
+ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13060__C1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ net1051 team_02_WB.instance_to_wrap.top.a1.row1\[121\] _03115_ _03290_ vssd1
+ vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15327_ clknet_leaf_45_wb_clk_i _01470_ _00140_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12539_ net347 net2155 net446 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14861__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15258_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[17\]
+ _00071_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14209_ net1256 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
X_15189_ net1142 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout408 _05809_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_2
XANTENNA__09582__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 net420 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_103_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] net758 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a22o_1
XANTENNA__09334__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09690__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ _04275_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or2_2
X_09681_ _05191_ _05193_ _05195_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__or4_1
X_08632_ net72 net1594 net957 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
XANTENNA__13416__S _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08563_ _03313_ _04171_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08494_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\] net979 vssd1 vssd1 vccd1
+ vccd1 _04190_ sky130_fd_sc_hd__or2_1
XANTENNA__10101__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout330_A _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1072_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\] net918 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\] net908 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\]
+ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_131_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout797_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13387__A net2477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11459__X _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10804__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10168__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
X_16779__1323 vssd1 vssd1 vccd1 vccd1 _16779__1323/HI net1323 sky130_fd_sc_hd__conb_1
Xhold495 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16698__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13106__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 _04515_ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08781__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_2
X_09948_ net514 _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__nor2_1
Xfanout942 _04532_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08768__X _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout953 _04455_ vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11117__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout964 net967 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_2
Xfanout975 _04284_ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_4
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XFILLER_0_204_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\] net781 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_129_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11910_ net236 net2189 net482 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
Xhold1162 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12230__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _05534_ _05537_ _07409_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__a21oi_1
Xhold1184 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_187_Left_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1195 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ net244 net2055 net493 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14560_ net1080 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
X_11772_ net240 net1954 net594 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XANTENNA__08944__A _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ team_02_WB.instance_to_wrap.top.pad.keyCode\[2\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__or4b_2
X_10723_ _06135_ _06239_ _06137_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_175_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ net1077 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_175_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16230_ clknet_leaf_6_wb_clk_i _02370_ _01038_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13442_ _02764_ _02763_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__nor2_1
XANTENNA_input93_A wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10654_ _06168_ _06170_ _06167_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a21o_2
XANTENNA__13042__C1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13593__B1 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16161_ clknet_leaf_104_wb_clk_i _02301_ _00969_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13373_ team_02_WB.instance_to_wrap.ramload\[2\] net1011 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[2\] sky130_fd_sc_hd__and2_1
X_10585_ net421 _06071_ net375 _06101_ _06086_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload18 clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_8
XANTENNA__08950__Y _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload29 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_8
XFILLER_0_180_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15112_ net1072 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XANTENNA__09775__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12324_ net295 net1872 net566 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16092_ clknet_leaf_16_wb_clk_i _02232_ _00900_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15043_ net1233 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
X_12255_ net290 net2088 net572 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12405__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11206_ net948 _06705_ _06711_ net607 vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__o211a_1
X_12186_ net271 net2186 net578 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15285__Q team_02_WB.instance_to_wrap.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08772__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11137_ _04951_ net664 _06643_ net795 _06644_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o221a_1
XANTENNA__09316__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ net371 _06510_ _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__o21ai_2
X_15945_ clknet_leaf_113_wb_clk_i _02085_ _00753_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] net791 net650 _05535_
+ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12140__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ clknet_leaf_36_wb_clk_i _02016_ _00684_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10331__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14827_ net1124 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14758_ net1213 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14689_ net1260 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
XANTENNA__11280__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ clknet_leaf_70_wb_clk_i net1418 _01236_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ clknet_leaf_39_wb_clk_i _02499_ _01167_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11279__X _06782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12315__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09555__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08763__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] net901 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a22o_1
Xfanout227 _03859_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07994_ _03692_ net256 _03686_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__a21oi_1
Xfanout249 _06498_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09307__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _05240_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout280_A _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10630__Y _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] net752 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a22o_1
XANTENNA__10322__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08615_ net80 net1442 net955 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09595_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] net816 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\]
+ _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08279__C1 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net1573 net792 net651 _04197_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08477_ _04175_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09794__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] net816 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\]
+ _05884_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09029_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\] net826 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\]
+ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12225__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ net350 net2222 net474 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__mux2_1
XANTENNA__09546__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 team_02_WB.instance_to_wrap.ramaddr\[11\] vssd1 vssd1 vccd1 vccd1 net1632
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08004__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold281 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 team_02_WB.instance_to_wrap.ramstore\[0\] vssd1 vssd1 vccd1 vccd1 net1654
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 _04376_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_4
Xfanout761 _04373_ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout772 _04371_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_195_Left_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991_ net1180 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_4
XANTENNA__11105__A2 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_4
XANTENNA__11365__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15730_ clknet_leaf_54_wb_clk_i _01870_ _00538_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12942_ team_02_WB.instance_to_wrap.top.pc\[20\] _06186_ vssd1 vssd1 vccd1 vccd1
+ _07462_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ clknet_leaf_49_wb_clk_i _01801_ _00469_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12873_ _07390_ _07392_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12066__A0 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14612_ net1241 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
X_11824_ net304 net2540 net589 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15592_ clknet_leaf_11_wb_clk_i _01732_ _00400_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10616__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14543_ net1222 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XANTENNA__10268__X _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ net308 net2166 net597 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10092__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _06222_ _06221_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and2b_1
X_14474_ net1188 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
X_11686_ _05966_ _07157_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__nand3_1
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16213_ clknet_leaf_31_wb_clk_i _02353_ _01021_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13425_ team_02_WB.instance_to_wrap.top.lcd.currentState\[3\] net962 vssd1 vssd1
+ vccd1 vccd1 _03035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__inv_2
Xclkload107 clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload107/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08680__Y _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__A1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16144_ clknet_leaf_30_wb_clk_i _02284_ _00952_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10568_ net424 net413 vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__nand2_1
XANTENNA__11041__B2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09785__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08613__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13356_ team_02_WB.instance_to_wrap.ramload\[18\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[18\] sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13318__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12307_ net352 net2218 net568 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12135__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16075_ clknet_leaf_17_wb_clk_i _02215_ _00883_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10444__A _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ _05986_ _05987_ _05989_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a22o_1
X_13287_ team_02_WB.instance_to_wrap.top.pc\[16\] net1054 _06807_ net933 vssd1 vssd1
+ vccd1 vccd1 _02993_ sky130_fd_sc_hd__a22o_1
X_15026_ net1258 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XANTENNA__09537__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ net1740 net360 net615 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_max_cap510_A _05533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ net332 net2260 net462 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13474__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15928_ clknet_leaf_121_wb_clk_i _02068_ _00736_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10304__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09170__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10855__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15859_ clknet_leaf_58_wb_clk_i _01999_ _00667_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08400_ _04102_ _04104_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__and3_1
XANTENNA__12057__A0 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _04890_ _04892_ _04894_ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__or4_1
X_08331_ _04024_ _04042_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16778__1322 vssd1 vssd1 vccd1 vccd1 _16778__1322/HI net1322 sky130_fd_sc_hd__conb_1
X_08262_ _03974_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__nand2_1
XANTENNA__10083__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08193_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03858_ vssd1 vssd1 vccd1
+ vccd1 _03911_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13649__B net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12045__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11884__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12965__A_N _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1202_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _03668_ _03699_ _03666_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10360__Y _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09716_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] net927 net809 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09161__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__A1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _05156_ _05160_ _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__or4_4
XFILLER_0_179_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout927_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09578_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\] net725 net717 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08529_ net1048 _04214_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13260__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ _05916_ _06003_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10074__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ net416 net665 _06536_ _06963_ net794 vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__o32a_1
XFILLER_0_162_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09216__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ net1491 net1020 net939 _04946_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a22o_1
X_10422_ _05292_ _05935_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_137_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14190_ net1075 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10353_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\] net753 net725 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13141_ net789 _07332_ _07510_ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13072_ _06623_ net234 _02848_ net978 _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o221a_1
XANTENNA__11079__B _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] net922 net804 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a22o_1
XANTENNA_input56_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net286 net2139 net475 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XANTENNA__11794__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13079__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _07209_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_6
Xfanout591 _07194_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_4
X_16762_ net1306 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
X_13974_ net1164 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_189_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15713_ clknet_leaf_103_wb_clk_i _01853_ _00521_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12925_ team_02_WB.instance_to_wrap.top.pc\[30\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _07445_ sky130_fd_sc_hd__nand2_1
X_16693_ clknet_leaf_70_wb_clk_i _02810_ _01417_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15644_ clknet_leaf_19_wb_clk_i _01784_ _00452_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12856_ _05314_ _06200_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__nand2_1
XANTENNA__08608__S _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11807_ net245 net2051 net589 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ clknet_leaf_120_wb_clk_i _01715_ _00383_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12787_ _06903_ _07308_ _07309_ _07310_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nor4_1
XANTENNA__11262__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14526_ net1130 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11738_ _04291_ net641 _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__or3_4
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11969__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10873__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14457_ net1091 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_11669_ _05271_ _05290_ _05990_ _07154_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] _03019_ vssd1 vssd1 vccd1
+ vccd1 _03020_ sky130_fd_sc_hd__nand2_1
XANTENNA__07748__A team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09758__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14388_ net1241 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08966__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ clknet_leaf_62_wb_clk_i _02267_ _00935_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13339_ team_02_WB.instance_to_wrap.ramload\[1\] net1018 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[1\] sky130_fd_sc_hd__and2_1
X_16058_ clknet_leaf_19_wb_clk_i _02198_ _00866_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11317__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07900_ _03521_ _03553_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15009_ net1135 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
X_08880_ net16 net1030 net987 net2520 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__o22a_1
XFILLER_0_209_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07831_ _03519_ _03552_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09930__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ _03481_ _03483_ _03484_ _03476_ _03461_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a32o_1
XANTENNA__09143__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] net911 net905 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a22o_1
X_07693_ _03384_ _03411_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ _04927_ _04947_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__nand2_1
XANTENNA__08518__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09363_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\] net728 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\]
+ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout243_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _04000_ _04018_ _04002_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10056__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11253__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] net912 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08245_ _03929_ _03959_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nand2_1
XANTENNA__11879__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1152_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__A team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _03852_ _03861_ _03889_ _03856_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09749__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08957__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout877_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__12503__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09382__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15957__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09134__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net382 _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ net848 _06161_ _06249_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__o31a_1
XFILLER_0_179_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10295__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13690_ net1139 _03215_ _03216_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ net245 net2050 net436 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10047__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ clknet_leaf_81_wb_clk_i _01500_ _00173_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_182_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12572_ net348 net2049 net443 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ net1173 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XANTENNA__11789__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11523_ net426 net385 _06297_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15291_ clknet_leaf_68_wb_clk_i _01435_ _00104_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08671__B team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ net1129 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
X_11454_ net668 _06937_ _06949_ net836 _06947_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_150_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10405_ _05919_ _05920_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nand2_1
X_14173_ net1181 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11385_ net954 _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13124_ _07375_ _07416_ _07374_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a21oi_1
X_10336_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] net796 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\]
+ _05852_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10267_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] net997 _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__a22o_1
X_13055_ team_02_WB.instance_to_wrap.top.pc\[26\] net1024 _02836_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01507_ sky130_fd_sc_hd__a22o_1
XANTENNA__12413__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16777__1321 vssd1 vssd1 vccd1 vccd1 _16777__1321/HI net1321 sky130_fd_sc_hd__conb_1
XANTENNA__09373__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ net352 net2567 net478 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XANTENNA__09912__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ net969 _05695_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_204_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16745_ net1290 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
X_13957_ net1249 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
XANTENNA__10286__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ _04971_ _06180_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o21ai_1
X_16676_ clknet_leaf_65_wb_clk_i _02793_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ net1250 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_196_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15627_ clknet_leaf_15_wb_clk_i _01767_ _00435_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12839_ _04802_ _06150_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15558_ clknet_leaf_6_wb_clk_i _01698_ _00366_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09979__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08100__B2 _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ net1120 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15489_ clknet_leaf_104_wb_clk_i _01629_ _00297_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08030_ net2461 net1007 net980 _03752_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13199__B _02953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput41 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
Xinput52 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xmax_cap500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_1
XFILLER_0_102_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold803 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_2
Xhold814 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08403__A2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold825 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput96 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
Xhold836 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09693__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold847 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold858 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\] net809 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08932_ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] net1010 _04232_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a221o_1
XANTENNA__12323__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10632__A team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ net150 net1040 net1037 net1417 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XANTENNA__08102__A team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07814_ _03499_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__xor2_2
XANTENNA__13943__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__X _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08794_ net548 _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or2_1
XANTENNA__09116__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07745_ _03461_ _03462_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1
+ vccd1 vccd1 _03468_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout458_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07678__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07676_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _03396_ _03397_ vssd1 vssd1
+ vccd1 vccd1 _03399_ sky130_fd_sc_hd__or3_1
X_09415_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] net913 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a22o_1
XANTENNA__08475__C team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10029__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ net533 _04861_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] net695 _04784_ _04787_
+ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08228_ _03943_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15378__Q team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11529__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08159_ _03865_ _03867_ _03876_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or3_1
X_11170_ _06672_ _06675_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__and3_1
XANTENNA__10201__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07602__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net905 net804 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\]
+ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12233__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13687__C1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09355__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\] net733 net713 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a22o_1
XANTENNA__13151__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ net1214 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
XANTENNA__16135__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ net1154 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__inv_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ net1180 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XANTENNA__08666__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16530_ clknet_leaf_82_wb_clk_i _00010_ _01337_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13742_ _03247_ _03248_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__nor2_1
XANTENNA__12662__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _04734_ _04778_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16461_ clknet_leaf_69_wb_clk_i net1606 _01269_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
X_13673_ net1527 _03206_ net1139 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a21oi_1
X_10885_ net391 _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__or2_1
XANTENNA__14684__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15412_ clknet_leaf_3_wb_clk_i _01552_ _00220_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ net1711 net298 net554 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__mux2_1
X_16392_ clknet_leaf_89_wb_clk_i _02527_ _01200_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15343_ clknet_leaf_73_wb_clk_i _01483_ _00156_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_12555_ net294 net1843 net444 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11506_ _06920_ _06998_ net396 vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__mux2_1
X_15274_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_read_i _00087_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.Ren sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ net289 net2326 net557 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14225_ net1229 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ team_02_WB.instance_to_wrap.top.pc\[11\] net973 _06933_ net1001 _06837_ vssd1
+ vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12932__A team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ net1216 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ _06014_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_210_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ net229 _02877_ _06786_ net232 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__inv_2
XANTENNA__10452__A _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ net1180 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
X_11299_ net379 _06571_ _06639_ _06567_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_165_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _06460_ net233 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nor2_1
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_4
XANTENNA__11982__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 net1170 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_2
XFILLER_0_178_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1172 net1175 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_4
Xfanout1183 net1187 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__buf_4
Xfanout1194 net1202 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_198_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13482__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09649__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14989_ net1160 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10259__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16728_ net1356 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_88_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16659_ clknet_leaf_93_wb_clk_i _02778_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09200_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] net915 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] net898 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a221o_1
XANTENNA__12318__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\] net723 _04577_ _04578_
+ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _03708_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__or2_1
Xhold600 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_116_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold622 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10633__Y _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12053__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\] net843 _05475_ _05477_
+ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a2111o_1
Xhold699 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1115_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ net1391 _04439_ net930 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
X_09895_ _05406_ _05408_ _05410_ _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__or4_1
XANTENNA__11144__B1 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11892__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_A _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11695__A1 _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ net148 net1039 net1037 net1508 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
X_08777_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\] net765 _04388_ _04393_
+ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout742_A _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07728_ _03445_ _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ _03353_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11480__X _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ net996 _05625_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12736__B _06851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16776__1320 vssd1 vssd1 vccd1 vccd1 _16776__1320/HI net1320 sky130_fd_sc_hd__conb_1
X_09329_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\] net864 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12228__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12340_ net350 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\] net564 vssd1
+ vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12271_ net358 net1915 net573 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ net1096 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11222_ net418 _06726_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09040__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _04997_ _06659_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09328__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] net778 _05617_ _05620_
+ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a211o_1
X_15961_ clknet_leaf_124_wb_clk_i _02101_ _00769_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11084_ net974 _06593_ _06592_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_147_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] net909 _05538_ _05551_
+ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__a211o_1
X_14912_ net1102 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
X_15892_ clknet_leaf_123_wb_clk_i _02032_ _00700_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08677__A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14843_ net1084 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11438__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14774_ net1106 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
X_11986_ net276 net2424 net478 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
X_16513_ clknet_leaf_0_wb_clk_i _02647_ _01320_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13725_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03017_ vssd1 vssd1 vccd1
+ vccd1 _03237_ sky130_fd_sc_hd__or2_1
X_10937_ net410 _06449_ _06359_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10110__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16444_ clknet_leaf_61_wb_clk_i net1435 _01252_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13656_ _04153_ net850 _03196_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a21oi_1
X_10868_ net367 _06055_ _06056_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__and3_1
XANTENNA__08616__S _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_183_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ net1805 net243 net554 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__mux2_1
X_16375_ clknet_leaf_87_wb_clk_i _02515_ _01183_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12138__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ team_02_WB.instance_to_wrap.top.a1.row2\[25\] _03118_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[105\]
+ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ net542 net387 _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15326_ clknet_leaf_71_wb_clk_i _01469_ _00139_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12538_ net351 net2537 net446 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11977__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15257_ clknet_leaf_106_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[16\]
+ _00070_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_12469_ net359 net1911 net452 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14208_ net1106 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XANTENNA__09567__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13477__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net1140 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10177__A1 _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09031__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ net1076 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
Xfanout409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_2
XANTENNA__09319__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13115__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ net1062 _04267_ net978 vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__o21ai_4
XANTENNA__13493__A _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\] net921 net901 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\]
+ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a221o_1
XANTENNA__12601__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ net83 net1548 net955 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04175_ vssd1 vssd1 vccd1
+ vccd1 _04231_ sky130_fd_sc_hd__or2_1
XANTENNA__09098__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ net1048 _04185_ _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a31o_1
XANTENNA__08845__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12837__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__X _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08526__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout323_A _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__inv_2
XANTENNA__11601__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09270__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09045_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] net900 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1232_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13387__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold441 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold474 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold485 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold496 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1118_X net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout910 _04523_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_4
Xfanout921 _04515_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
Xfanout932 _04335_ vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
X_09947_ _05444_ net623 net968 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__mux2_2
Xfanout943 _04532_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout954 _04455_ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout957_A _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_2
Xfanout976 net977 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12511__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\] net745 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a22o_1
Xfanout987 _04432_ vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 _04264_ vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15698__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1130 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09730__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1152 team_02_WB.instance_to_wrap.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net2514
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ net1605 net1041 net991 team_02_WB.instance_to_wrap.ramaddr\[2\] vssd1 vssd1
+ vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
Xhold1163 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1174 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1196 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net242 net2549 net492 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XANTENNA__09089__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11771_ _04291_ _04333_ net642 _06280_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__or4_4
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13290__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__B _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13510_ net1505 net1363 _03071_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__mux2_1
X_10722_ team_02_WB.instance_to_wrap.top.pc\[28\] _06140_ _06238_ vssd1 vssd1 vccd1
+ vccd1 _06239_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14490_ net1089 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ net1067 _03028_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ team_02_WB.instance_to_wrap.top.a1.instruction\[24\] _04283_ _06169_ vssd1
+ vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16160_ clknet_leaf_109_wb_clk_i _02300_ _00968_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11053__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input86_A wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13372_ net1601 net1012 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ _06093_ _06100_ net397 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload19 clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11797__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15111_ net1113 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net286 net1791 net567 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16091_ clknet_leaf_34_wb_clk_i _02231_ _00899_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09549__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ net1230 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
X_12254_ net276 net2102 net572 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11205_ _04284_ _06710_ _06709_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_71_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12185_ net263 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] net578 vssd1
+ vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ _04948_ net661 net658 _04949_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__a22oi_1
X_11067_ net371 _06576_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__nand2_1
XANTENNA__12421__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15944_ clknet_leaf_24_wb_clk_i _02084_ _00752_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09721__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10018_ _04421_ _05441_ net550 vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15875_ clknet_leaf_27_wb_clk_i _02015_ _00683_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14826_ net1127 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14757_ net1173 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
X_11969_ net359 net2468 net587 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13708_ net2201 _03226_ net1066 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14688_ net1105 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11280__B _06782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ net1500 net963 _03187_ _00018_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__o211a_1
X_16427_ clknet_leaf_83_wb_clk_i net1504 _01235_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ clknet_leaf_7_wb_clk_i _02498_ _01166_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09252__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15309_ clknet_leaf_72_wb_clk_i _01452_ _00122_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16289_ clknet_leaf_101_wb_clk_i _02429_ _01097_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10624__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09972__Y _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09801_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\] net810 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__a221o_1
XANTENNA__09960__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15840__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07993_ _03686_ _03692_ net256 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__and3_1
Xfanout239 _06424_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
X_09732_ _05242_ _05244_ _05246_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or4_2
XANTENNA__12331__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\] net771 _05170_ _05173_
+ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a2111o_1
X_08614_ net81 net1535 net955 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13951__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1019_A team_02_WB.instance_to_wrap.ramload\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09594_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] net926 net906 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ net2451 net792 net651 _04194_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XANTENNA__13272__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08476_ _04169_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09491__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10087__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13024__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14782__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09779__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire629 _05121_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12573__Y _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12506__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\] net915 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 team_02_WB.instance_to_wrap.top.a1.row2\[9\] vssd1 vssd1 vccd1 vccd1 net1622
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_02_WB.instance_to_wrap.ramaddr\[18\] vssd1 vssd1 vccd1 vccd1 net1633
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 team_02_WB.instance_to_wrap.top.a1.row1\[0\] vssd1 vssd1 vccd1 vccd1 net1655
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 _04379_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_4
Xfanout751 _04376_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12241__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout762 _04373_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13990_ net1212 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XANTENNA__10550__A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout773 _04369_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_8
Xfanout784 _04366_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
Xfanout795 _06105_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09703__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ team_02_WB.instance_to_wrap.top.pc\[20\] _06186_ vssd1 vssd1 vccd1 vccd1
+ _07461_ sky130_fd_sc_hd__nor2_1
X_15660_ clknet_leaf_2_wb_clk_i _01800_ _00468_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12872_ _07389_ _07391_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_177_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14611_ net1079 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ net296 net1939 net590 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__mux2_1
X_15591_ clknet_leaf_41_wb_clk_i _01731_ _00399_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14542_ net1075 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
X_11754_ net302 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\] net598 vssd1
+ vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10705_ team_02_WB.instance_to_wrap.top.pc\[19\] _06186_ vssd1 vssd1 vccd1 vccd1
+ _06222_ sky130_fd_sc_hd__xnor2_1
X_14473_ net1216 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ net542 _04692_ _05967_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16212_ clknet_leaf_3_wb_clk_i _02352_ _01020_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13424_ _03030_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10636_ _04344_ _04349_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_155_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08690__A _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09234__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload108 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__inv_8
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12924__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16143_ clknet_leaf_43_wb_clk_i _02283_ _00951_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11041__A2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ net1552 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[17\]
+ sky130_fd_sc_hd__and2_1
X_10567_ net420 net409 vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__nor2_1
XANTENNA__12416__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ net365 net2231 net568 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16074_ clknet_leaf_32_wb_clk_i _02214_ _00882_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13286_ net1629 net984 net966 _02992_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_188_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10498_ _05991_ _06013_ _05990_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__o21a_1
X_15025_ net1233 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
X_12237_ net2238 net342 net613 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08689__X _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ net336 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\] net465 vssd1
+ vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
X_11119_ _04951_ _05947_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_207_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12151__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ net1653 net327 net581 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_X clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15927_ clknet_leaf_120_wb_clk_i _02067_ _00735_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11990__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ clknet_leaf_54_wb_clk_i _01998_ _00666_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809_ net1088 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15789_ clknet_leaf_49_wb_clk_i _01929_ _00597_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10068__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ _04024_ _04035_ _04040_ _04039_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__Y _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08261_ _03952_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08192_ _03872_ _03896_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09225__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12834__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12326__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14107__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13309__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13946__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_A _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09933__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _03660_ _03664_ _03673_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__o21ba_1
X_09715_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] net889 net863 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout655_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09646_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] net900 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\]
+ _05147_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a221o_1
XANTENNA__10846__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_182_Right_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09577_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\] net769 net685 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout822_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08528_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\] net979 vssd1 vssd1 vccd1
+ vccd1 _04215_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09464__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08459_ _03307_ _04154_ _04160_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11470_ net376 _06773_ _06961_ net382 _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09216__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11559__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10421_ _05292_ _05936_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10545__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12236__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08975__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ _07479_ _07481_ _07509_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__nor3_1
XANTENNA__10231__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10352_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] net757 _05858_ _05861_
+ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_20_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07632__D1 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ net231 _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__nand2_1
XANTENNA__12760__A _04694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10283_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] net940 _05796_ _05797_
+ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13180__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ net272 net2094 net476 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
XANTENNA_input49_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_X clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15266__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_4
Xfanout581 _07209_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_4
Xfanout592 net593 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13195__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16761_ net1305 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_45_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13973_ net1160 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XFILLER_0_205_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10298__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15712_ clknet_leaf_109_wb_clk_i _01852_ _00520_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12924_ team_02_WB.instance_to_wrap.top.pc\[30\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _07444_ sky130_fd_sc_hd__or2_1
X_16692_ clknet_leaf_70_wb_clk_i _02809_ _01416_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08685__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09133__X _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15643_ clknet_leaf_33_wb_clk_i _01783_ _00451_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _05314_ _06200_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11806_ net243 net2090 net589 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
X_15574_ clknet_leaf_21_wb_clk_i _01714_ _00382_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12786_ _06722_ _06753_ _06770_ _06802_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09455__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14525_ net1181 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11737_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__or3b_4
XANTENNA__11262__A2 _06759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13133__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14456_ net1195 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
X_11668_ _05993_ _07152_ _07153_ _05991_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_54_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09207__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13407_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__and2_1
X_10619_ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12146__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ net1078 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
X_11599_ net2046 net357 net640 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16126_ clknet_leaf_4_wb_clk_i _02266_ _00934_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13338_ net2397 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[0\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11985__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16057_ clknet_leaf_125_wb_clk_i _02197_ _00865_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13269_ team_02_WB.instance_to_wrap.top.pc\[25\] net1055 net934 _02983_ vssd1 vssd1
+ vccd1 vccd1 _02984_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15008_ net1160 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XANTENNA__09915__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07830_ _03511_ _03519_ _03534_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__or3_1
XANTENNA__09027__Y _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire623_A _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ _03453_ _03463_ _03480_ _03448_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a22o_1
XANTENNA__15759__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14597__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07692_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__inv_2
X_09431_ _04927_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\] net764 net736 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09446__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08313_ _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__or2_1
XANTENNA__11253__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\] net814 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ _04807_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_72_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12845__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net2429 net1007 net980 _03960_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XANTENNA__08534__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12056__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _03888_ _03862_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__nand2b_1
XANTENNA_clkbuf_4_6__f_wb_clk_i_X clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1145_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11895__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__15289__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09906__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07674__A team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__B2 _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_81_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1100_X net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _03652_ _03655_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ net400 _06106_ _06480_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_168_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09685__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09629_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\] net727 _05141_ _05142_
+ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a2111oi_2
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ net243 net2133 net436 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input103_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ net352 net2099 net442 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__mux2_1
XANTENNA__08645__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14310_ net1204 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11522_ _05649_ _06004_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15290_ clknet_leaf_70_wb_clk_i _01434_ _00103_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08671__C team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ net1260 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16064__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11453_ _05927_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10204__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ _05579_ _05603_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07605__D1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14172_ net1201 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
X_11384_ net668 _06867_ _06882_ net836 _06880_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__o221a_1
XFILLER_0_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13123_ _07513_ _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_185_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10335_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] net926 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ net977 _07435_ _02834_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__o31ai_1
X_10266_ _05763_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__nand2_1
X_12005_ net363 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\] net478 vssd1
+ vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
X_10197_ net971 net620 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_204_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16744_ net1289 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__08619__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ net1240 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XANTENNA__09676__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12907_ _07365_ _07367_ _07425_ _06184_ _05017_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__a32o_1
X_16675_ clknet_leaf_65_wb_clk_i _02792_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11483__A2 _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887_ net1246 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XFILLER_0_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15626_ clknet_leaf_37_wb_clk_i _01766_ _00434_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12838_ net539 _06147_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_196_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09428__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ net663 _07177_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__o21ai_1
X_15557_ clknet_leaf_28_wb_clk_i _01697_ _00365_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14508_ net1209 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12983__A2 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15488_ clknet_leaf_18_wb_clk_i _01628_ _00296_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ net1182 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_2
Xinput53 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09061__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput75 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold804 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
Xhold826 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09600__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_2
Xinput97 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_92_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold837 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ clknet_leaf_49_wb_clk_i _02249_ _00917_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold848 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12604__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] net917 net907 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a22o_1
Xhold859 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] net959 _04221_ _04173_ vssd1
+ vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08862_ net161 net1046 net1037 net1501 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11171__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _03532_ _03533_ _03502_ _03510_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a211o_1
X_08793_ net650 _04420_ _04421_ net791 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__a22oi_4
X_07744_ _03435_ _03463_ _03464_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11459__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07675_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or2_1
XANTENNA__08875__B1 _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09414_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] net928 net811 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1095_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09419__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ _04842_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1262_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\] net758 _04789_ _04790_
+ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08227_ _03909_ _03915_ _03926_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__or3_1
XANTENNA__14790__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08158_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout987_A _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07602__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10823__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ _03755_ _03786_ _03782_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o21a_2
XANTENNA__12514__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] net910 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] net765 net737 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a22o_1
XANTENNA__13151__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ net1154 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__inv_2
X_14790_ net1213 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09658__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ net2587 _03245_ net951 vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_119_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10953_ net1591 net253 net639 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08866__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11941__X _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10673__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ _03202_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] _03200_ _03205_
+ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__or4bb_2
X_16460_ clknet_leaf_84_wb_clk_i net1575 _01268_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_10884_ _06080_ _06081_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15411_ clknet_leaf_47_wb_clk_i _01551_ _00219_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12623_ net2109 net308 net555 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16391_ clknet_leaf_89_wb_clk_i _02526_ _01199_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ clknet_leaf_84_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] _00155_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[3\] sky130_fd_sc_hd__dfrtp_1
X_12554_ net287 net2580 net443 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XANTENNA__09291__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _06959_ _06997_ net367 vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__mux2_1
X_15273_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_write_i _00086_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.Wen sky130_fd_sc_hd__dfrtp_2
X_12485_ net276 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] net556 vssd1
+ vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__mux2_1
X_14224_ net1258 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11436_ _06259_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_128_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09043__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12932__B _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14155_ net1124 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XANTENNA__12424__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ _05377_ _06013_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10292__X _05809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ _07369_ _07370_ _07421_ net976 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a31o_1
X_10318_ net791 _05442_ _05834_ _04331_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__a22oi_4
X_14086_ net1212 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
X_11298_ _05207_ net660 net657 _05210_ _06799_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a221o_1
XANTENNA__13678__B1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _02821_ _02818_ _07349_ team_02_WB.instance_to_wrap.top.pc\[29\] vssd1 vssd1
+ vccd1 vccd1 _01510_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_119_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10249_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] net703 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_4
XANTENNA__09897__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_2
Xfanout1162 net1163 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_4
XFILLER_0_206_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10900__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1173 net1175 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net1187 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_198_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11564__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1195 net1198 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
XFILLER_0_89_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09649__A2 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14988_ net1154 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16727_ net1355 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XANTENNA__08857__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ net1164 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16658_ clknet_leaf_94_wb_clk_i _02777_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08609__A0 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15609_ clknet_leaf_125_wb_clk_i _01749_ _00417_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16589_ clknet_leaf_90_wb_clk_i _02708_ _01382_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] net804 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__a22o_1
XANTENNA__09282__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09061_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\] net715 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ _03694_ net256 _03680_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09034__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__A1 team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold612 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__B _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 team_02_WB.instance_to_wrap.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net1996
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12334__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold645 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold656 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold667 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\] net786 _05478_ _05479_
+ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a211o_1
Xhold689 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ net1047 _04203_ _04214_ net1009 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a32o_1
XANTENNA__13954__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\] net870 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ _05403_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__a221o_1
XANTENNA__09888__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08845_ net149 net1043 net1035 net1415 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout470_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__Y _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\] net781 _04396_ _04398_
+ _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a2111o_1
X_07727_ _03410_ net425 _03415_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08848__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14785__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03349_ vssd1 vssd1 vccd1
+ vccd1 _03381_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12509__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ team_02_WB.instance_to_wrap.top.a1.state\[2\] _03313_ vssd1 vssd1 vccd1 vccd1
+ _03314_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout902_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1265_X net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09328_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] net916 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08076__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09273__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09259_ net971 _04774_ net544 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_173_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12270_ net344 net1751 net574 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ net413 _06483_ _06717_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11649__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13235__B1_N net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12244__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _05042_ _06600_ _05039_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__o21a_1
XANTENNA__08023__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10103_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\] net748 _05618_ _05619_
+ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a211o_1
X_15960_ clknet_leaf_121_wb_clk_i _02100_ _00768_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11083_ _06173_ _06231_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09879__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10034_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] net892 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\]
+ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__a221o_1
X_14911_ net1108 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
X_15891_ clknet_leaf_58_wb_clk_i _02031_ _00699_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14842_ net1096 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11438__A2 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ net281 net2220 net479 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
X_14773_ net1200 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16512_ clknet_leaf_127_wb_clk_i _02646_ _01319_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ net410 _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__nor2_1
X_13724_ _03018_ net950 _03236_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16443_ clknet_leaf_61_wb_clk_i net1488 _01251_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
X_10867_ _06378_ _06380_ net395 vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__mux2_1
X_13655_ net1385 net850 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__nor2_1
XANTENNA__12419__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10728__A _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12606_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] net642 _06277_ _06279_
+ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13586_ team_02_WB.instance_to_wrap.top.a1.row1\[113\] _03121_ _03124_ team_02_WB.instance_to_wrap.top.a1.row2\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a22o_1
XANTENNA__08980__X _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13060__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16374_ clknet_leaf_21_wb_clk_i _02514_ _01182_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10798_ _04714_ net387 vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13060__B2 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15325_ clknet_leaf_61_wb_clk_i _01468_ _00138_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11071__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ net364 net2183 net446 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08632__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15256_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[15\]
+ _00069_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_12468_ net342 net1840 net451 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _06011_ net663 vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__nor2_1
X_14207_ net1115 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XANTENNA__12154__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ net1140 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
X_12399_ net336 net2284 net461 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ net1090 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XANTENNA__11993__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13115__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ net1257 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XANTENNA_wire536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ net94 net1624 net956 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04175_ vssd1 vssd1 vccd1
+ vccd1 _04230_ sky130_fd_sc_hd__nor2_1
X_08492_ team_02_WB.instance_to_wrap.top.a1.row1\[19\] net849 vssd1 vssd1 vccd1 vccd1
+ _04189_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10101__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12837__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12329__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ _04623_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor2_8
XANTENNA__13949__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12853__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1058_A team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13301__X _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\] net891 _04551_ _04560_
+ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1166_A team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12064__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12562__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10168__A2 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 _04526_ vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_8
Xfanout911 _04523_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_4
Xhold497 team_02_WB.instance_to_wrap.top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net1859
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08781__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout922 _04513_ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_4
X_09946_ _05456_ _05459_ _05461_ _05462_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__nor4_2
XANTENNA__11117__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout933 net935 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
Xfanout944 _04501_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_2
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_2
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
Xhold1120 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\] net689 _05382_ _05393_
+ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_2
Xhold1142 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ net131 net1045 net992 net1429 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
Xhold1153 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\] net713 net705 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1197 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ net346 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] net596 vssd1
+ vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
XANTENNA__09494__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13290__B2 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ _06145_ _06237_ _06141_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__o21a_1
XANTENNA__10548__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _03034_ _03041_ _03042_ _03045_ _03046_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a32o_1
X_10652_ net996 _04492_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__or2_1
XANTENNA__09246__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13042__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13042__B2 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13371_ net2397 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[0\]
+ sky130_fd_sc_hd__and2_1
X_10583_ _06096_ _06099_ net373 vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ net272 net2464 net565 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__mux2_1
X_15110_ net1074 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16090_ clknet_leaf_50_wb_clk_i _02230_ _00898_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input79_A wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15041_ net1245 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
X_12253_ net283 net2056 net573 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XANTENNA__10159__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11204_ _06224_ _06225_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12184_ net265 net2004 net578 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ net423 _06634_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__nand2_1
XANTENNA__08772__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12702__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12305__A0 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11108__B2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_196_Right_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13648__A3 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__A team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11066_ _06321_ _06324_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__nor2_1
X_15943_ clknet_leaf_40_wb_clk_i _02083_ _00751_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ net509 vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15874_ clknet_leaf_119_wb_clk_i _02014_ _00682_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10331__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14825_ net1210 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12938__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_176_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15792__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14756_ net1092 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
XANTENNA__09485__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13281__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ net343 net1742 net585 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13707_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] _03226_ vssd1 vssd1 vccd1
+ vccd1 _03227_ sky130_fd_sc_hd__and2_1
X_10919_ _06293_ _06299_ net367 vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12149__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14687_ net1116 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_11899_ net340 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] net489 vssd1
+ vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux2_1
X_16426_ clknet_leaf_82_wb_clk_i _02561_ _01234_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ _03109_ _03113_ _03117_ team_02_WB.instance_to_wrap.top.a1.row1\[60\] _03023_
+ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11988__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16357_ clknet_leaf_28_wb_clk_i _02497_ _01165_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13569_ net1050 net1052 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03103_
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__and4_1
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12792__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15308_ clknet_leaf_82_wb_clk_i _01451_ _00121_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16288_ clknet_leaf_109_wb_clk_i _02428_ _01096_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15239_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[30\]
+ _00052_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_113_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] net916 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__a22o_1
XANTENNA__08763__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12612__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07992_ _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__nand2_1
Xfanout229 _07333_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09731_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\] net825 net873 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\]
+ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a221o_1
XANTENNA_wire539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\] net845 _05175_ _05176_
+ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10322__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ net82 net1534 net956 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
X_09593_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\] net796 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\]
+ _05105_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a221o_1
XANTENNA__10973__A2_N net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ net1599 net792 net651 _04191_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10086__A1 _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 _04174_
+ sky130_fd_sc_hd__nand3b_1
XANTENNA_fanout433_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12059__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1175_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11898__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire608 _05781_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_2
XFILLER_0_135_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire619 _05806_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_4
XANTENNA__13285__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout600_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09027_ _04516_ _04527_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11338__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold250 team_02_WB.instance_to_wrap.ramaddr\[24\] vssd1 vssd1 vccd1 vccd1 net1612
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09400__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 team_02_WB.instance_to_wrap.ramload\[31\] vssd1 vssd1 vccd1 vccd1 net1623
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 team_02_WB.instance_to_wrap.ramaddr\[25\] vssd1 vssd1 vccd1 vccd1 net1634
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_02_WB.instance_to_wrap.top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 net1645
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12522__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net732 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_6
Xfanout741 _04378_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_4
XANTENNA__16498__Q team_02_WB.START_ADDR_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08939__C _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout752 _04376_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
X_09929_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\] net824 net820 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout763 _04373_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout774 _04369_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_4
Xfanout796 net799 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_8
X_12940_ team_02_WB.instance_to_wrap.top.pc\[21\] _06184_ vssd1 vssd1 vccd1 vccd1
+ _07460_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11510__B2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ _05788_ net498 vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_177_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ net1185 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11822_ net308 net1526 net591 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XANTENNA__09467__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ clknet_leaf_8_wb_clk_i _01730_ _00398_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13263__B2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11274__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ net1122 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11753_ net295 net1493 net598 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ team_02_WB.instance_to_wrap.top.pc\[18\] _06188_ _06220_ vssd1 vssd1 vccd1
+ vccd1 _06221_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _04781_ _05968_ _05969_ _06373_ _07158_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09219__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14472_ net1111 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ clknet_leaf_51_wb_clk_i _02351_ _01019_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13423_ net1066 _03028_ _03031_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and3_1
X_10635_ team_02_WB.instance_to_wrap.top.pc\[25\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _06152_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11577__A1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload109/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ clknet_leaf_47_wb_clk_i _02282_ _00950_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13354_ net2631 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[16\]
+ sky130_fd_sc_hd__and2_1
X_10566_ net373 _06079_ _06080_ _06082_ net396 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12305_ net357 net2382 net570 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__mux2_1
XANTENNA__13318__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16073_ clknet_leaf_113_wb_clk_i _02213_ _00881_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13285_ _06782_ _02959_ team_02_WB.instance_to_wrap.top.pc\[17\] net1054 vssd1 vssd1
+ vccd1 vccd1 _02992_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11329__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10497_ _05336_ _05932_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_188_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15024_ net1258 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
X_12236_ net2142 net340 net613 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12432__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ net327 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\] net463 vssd1
+ vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ net1723 net271 net639 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
X_12098_ net1643 net322 net580 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _06268_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or2_1
X_15926_ clknet_leaf_22_wb_clk_i _02066_ _00734_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10304__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_188_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09170__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ clknet_leaf_128_wb_clk_i _01997_ _00665_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15044__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14808_ net1196 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XANTENNA__09458__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15788_ clknet_leaf_2_wb_clk_i _01928_ _00596_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14739_ net1073 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08260_ _03925_ _03960_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16409_ clknet_leaf_100_wb_clk_i _02544_ _01217_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_08191_ _03868_ _03905_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_99_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12607__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09630__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10635__B _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13309__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08599__Y _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10651__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09217__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _03684_ _03693_ _03697_ _03680_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09714_ net610 vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09697__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09161__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09645_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\] net834 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\]
+ _05161_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09576_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\] net838 _05090_ _05092_
+ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a211o_1
XFILLER_0_210_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ team_02_WB.instance_to_wrap.top.a1.data\[2\] net959 vssd1 vssd1 vccd1 vccd1
+ _04214_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout815_A _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ net1597 net1006 net981 _04161_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_172_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11008__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12517__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08389_ _04094_ _04096_ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10420_ _05936_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__inv_2
XANTENNA__11559__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09621__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] net777 _05862_ _05864_
+ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07632__C1 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__A2 _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _07457_ _07527_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10282_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\] net812 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\]
+ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net289 net1726 net475 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout560 net563 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_6
XFILLER_0_205_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout571 _07217_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_4
X_16760_ net1304 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
Xfanout582 _07209_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_6
Xfanout593 _07192_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_4
X_13972_ net1160 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
X_15711_ clknet_leaf_59_wb_clk_i _01851_ _00519_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09152__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12923_ _07441_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__xnor2_1
X_16691_ clknet_leaf_70_wb_clk_i _02808_ _01415_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08685__B team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15642_ clknet_leaf_50_wb_clk_i _01782_ _00450_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ net609 _06197_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_202_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ _04292_ net641 _07193_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__or3_1
X_15573_ clknet_leaf_31_wb_clk_i _01713_ _00381_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12785_ _06070_ _06313_ _06388_ net422 vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__o31a_1
XFILLER_0_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08972__Y _04489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09797__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524_ net1199 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
X_11736_ net348 net2386 net600 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08905__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15830__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10470__A1 _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14455_ net1210 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XANTENNA__12427__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ _05440_ _05464_ _05992_ _05376_ _05356_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__o32a_1
XFILLER_0_154_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13406_ _03300_ _03016_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10618_ team_02_WB.instance_to_wrap.top.pc\[29\] _06134_ vssd1 vssd1 vccd1 vccd1
+ _06135_ sky130_fd_sc_hd__nand2_1
XANTENNA__08206__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ net947 _07083_ _07086_ net605 vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__o211a_1
X_14386_ net1183 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
X_16125_ clknet_leaf_10_wb_clk_i _02265_ _00933_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08966__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10549_ _06064_ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10222__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13337_ net1057 team_02_WB.instance_to_wrap.top.ru.state\[2\] vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_iready sky130_fd_sc_hd__and2b_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16056_ clknet_leaf_114_wb_clk_i _02196_ _00864_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13268_ _06556_ _06588_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_209_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15007_ net1135 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
X_12219_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\] net270 net614 vssd1
+ vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__mux2_1
XANTENNA__12162__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ net1019 _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__nor2_4
XFILLER_0_209_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ _03457_ _03475_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__xor2_4
XANTENNA__09679__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13475__A1 team_02_WB.START_ADDR_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ clknet_leaf_28_wb_clk_i _02049_ _00717_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_07691_ _03372_ _03405_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_108_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08595__B net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09430_ net969 _04946_ _04497_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\] net747 _04867_ _04870_
+ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_121_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08312_ _03997_ _04018_ _03999_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\] net818 net908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\]
+ _04806_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09851__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _03932_ _03959_ _03929_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_103_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09500__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12337__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14118__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ _03892_ _03889_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__nand2b_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09603__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13957__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12861__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1040_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout598_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__clkbuf_4
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__12072__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA__09382__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _03657_ _03678_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_199_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09134__A2 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03609_ _03610_ vssd1 vssd1
+ vccd1 vccd1 _03612_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\] net746 _05143_ _05144_
+ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] net913 net885 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\]
+ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_194_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12570_ net364 net2247 net442 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09842__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11521_ net1542 net331 net637 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12247__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10556__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11452_ _05468_ _05926_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__nor2_1
X_14240_ net1102 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XANTENNA__08671__D team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire235 _07326_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_152_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10403_ net506 _05603_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__or2_1
X_14171_ net1087 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XANTENNA__07605__C1 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11383_ _06014_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12771__A _06942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15233__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\] net824 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a221o_1
XANTENNA_input61_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _07471_ _07472_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_185_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ net230 _02833_ _06526_ net233 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_76_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ net608 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__inv_2
X_12004_ net355 net1770 net480 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09373__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _05706_ _05709_ _05710_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nor4_2
XANTENNA__15383__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout390 net392 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
XFILLER_0_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09125__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16743_ net1288 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13955_ net1240 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12906_ _07367_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__nand2_1
X_16674_ clknet_leaf_65_wb_clk_i _02791_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13209__B2 _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10140__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ net1167 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
X_15625_ clknet_leaf_116_wb_clk_i _01765_ _00433_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_196_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ _04714_ _06143_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15556_ clknet_leaf_35_wb_clk_i _01696_ _00364_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12768_ _07277_ _07280_ _07281_ _07291_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__o22a_1
XANTENNA__09833__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14507_ net1098 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XANTENNA__12157__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11719_ net292 net1687 net600 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
X_15487_ clknet_leaf_62_wb_clk_i _01627_ _00295_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12699_ net344 net2198 net431 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14438_ net1213 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_1
XFILLER_0_140_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
XFILLER_0_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11996__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput43 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput54 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
X_14369_ net1256 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold805 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xinput65 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
Xhold816 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap524 net525 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_2
Xinput76 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput87 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_1
X_16108_ clknet_leaf_2_wb_clk_i _02248_ _00916_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold827 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xinput98 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
Xhold838 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13145__B1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16039_ clknet_leaf_39_wb_clk_i _02179_ _00847_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_08930_ net1406 _04449_ _04433_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ net1459 net1044 net1036 team_02_WB.instance_to_wrap.ramstore\[3\] vssd1 vssd1
+ vccd1 vccd1 _02565_ sky130_fd_sc_hd__a22o_1
X_07812_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__nand2_1
XANTENNA__12620__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] _04330_ net649 team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a22o_1
XANTENNA__09116__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03398_ _03432_ vssd1 vssd1
+ vccd1 vccd1 _03466_ sky130_fd_sc_hd__or3_1
XANTENNA_wire619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _03393_ _03394_ vssd1 vssd1
+ vccd1 vccd1 _03397_ sky130_fd_sc_hd__and3_1
XANTENNA__08875__A1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] net896 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12856__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1088_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ net970 net633 net543 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__o21a_1
XANTENNA__08627__A1 team_02_WB.START_ADDR_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_205_Left_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09275_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\] net844 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\]
+ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a221o_1
XANTENNA__12067__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1255_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ _03905_ _03914_ _03927_ _03908_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_43_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _03872_ _03873_ _03874_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__or3_2
XFILLER_0_133_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1043_X net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08088_ _03801_ _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__or2_1
XANTENNA__07602__A2 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09355__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\] net842 net681 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\]
+ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12530__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13740_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] _03245_ vssd1 vssd1 vccd1
+ vccd1 _03247_ sky130_fd_sc_hd__and2_1
XANTENNA__10122__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ net946 _06458_ _06465_ net605 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__o211a_2
XFILLER_0_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13671_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03201_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__and4bb_1
X_10883_ _06392_ _06393_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__o21a_1
XANTENNA__15142__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15410_ clknet_leaf_54_wb_clk_i _01550_ _00218_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12622_ net1897 net302 net553 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__mux2_1
XANTENNA__09411__Y _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16390_ clknet_leaf_89_wb_clk_i _02525_ _01198_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15341_ clknet_leaf_85_wb_clk_i _00009_ _00154_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ net275 net1847 net444 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XANTENNA__14981__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ _06049_ _06055_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__nand2b_1
XANTENNA__16181__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15272_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[31\]
+ _00085_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_12484_ net280 net2558 net558 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14223_ net1220 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
X_11435_ team_02_WB.instance_to_wrap.top.pc\[11\] _06258_ vssd1 vssd1 vccd1 vccd1
+ _06932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07595__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14154_ net1118 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
X_11366_ net1795 net296 net640 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10317_ _05785_ _04419_ net550 vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__mux2_1
X_13105_ _07369_ _07370_ _07421_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a21oi_1
X_11297_ _05211_ _06111_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__nor2_1
X_14085_ net1172 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
XANTENNA__15899__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10248_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\] net754 net751 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a22o_1
X_13036_ _06422_ net233 _02820_ net977 _07337_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__o221a_1
XFILLER_0_206_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1130 net1131 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_4
Xfanout1141 net1146 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_2
X_10179_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] net896 net943 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a22o_1
XANTENNA__12440__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1152 net1170 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_2
Xfanout1163 net1169 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__buf_4
Xfanout1174 net1175 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_2
XFILLER_0_206_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_4
XFILLER_0_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_198_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1196 net1198 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_4
X_14987_ net1135 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16726_ net1354 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13938_ net1229 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10113__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11861__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16657_ clknet_leaf_94_wb_clk_i _02776_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13869_ net1163 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
X_15608_ clknet_leaf_121_wb_clk_i _01748_ _00416_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09806__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16588_ clknet_leaf_92_wb_clk_i _02707_ _01381_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09050__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15539_ clknet_leaf_57_wb_clk_i _01679_ _00347_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11613__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14891__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09060_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] net775 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _03681_ _03713_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__xor2_2
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11579__X _07069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12615__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold602 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__A2 _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09585__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold635 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload33_A clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\] net750 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09337__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ net1409 _04438_ net930 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
X_09893_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] net820 net816 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\]
+ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout296_A _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12350__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ net1465 net1039 net1037 team_02_WB.instance_to_wrap.ramstore\[20\] vssd1
+ vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
X_08775_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] net681 net838 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\]
+ _04401_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a221o_1
XANTENNA__16054__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_A _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07726_ _03406_ _03438_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__xor2_2
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07657_ _03345_ _03347_ _03351_ _03361_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout728_A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07588_ team_02_WB.instance_to_wrap.top.a1.state\[1\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nor2_1
X_09327_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] net818 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__a22o_1
XANTENNA__12736__D _06901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08076__A2 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09258_ net971 _04774_ net544 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__o21a_1
X_08209_ _03897_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a21o_2
X_09189_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\] net735 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\]
+ _04705_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a221o_1
XANTENNA__12525__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10834__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_177_Right_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11220_ _05974_ net664 _06723_ net666 _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09576__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _04997_ _05946_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09119__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__B team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10102_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\] net786 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a22o_1
XANTENNA__09328__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11082_ net999 _06590_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__o21ba_1
X_10033_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] net823 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__a22o_1
X_14910_ net1188 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
XANTENNA__12260__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ clknet_leaf_76_wb_clk_i _02030_ _00698_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10343__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__A1 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ net1100 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ net1238 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11984_ _06626_ net2176 net479 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XANTENNA__08974__A team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16511_ clknet_leaf_127_wb_clk_i _02645_ _01318_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13723_ _03300_ _03016_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__nand2_1
X_10935_ net407 _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16442_ clknet_leaf_42_wb_clk_i net1413 _01250_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_193_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ net1380 _04161_ net850 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10866_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12605_ net346 net2366 net438 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16373_ clknet_leaf_31_wb_clk_i _02513_ _01181_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13585_ net1438 net962 _03139_ net1067 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__o211a_1
X_10797_ _06296_ _06312_ net412 vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15324_ clknet_leaf_45_wb_clk_i _01467_ _00137_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ net356 net1690 net448 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
XANTENNA__08913__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15255_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[14\]
+ _00068_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07596__Y _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ net338 net2171 net451 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__mux2_1
XANTENNA__12435__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13024__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ net1127 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _06010_ _06011_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09567__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15186_ net1140 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12398_ net327 net2313 net459 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__mux2_1
XANTENNA__08775__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ net1090 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
X_11349_ _06745_ _06848_ net397 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09319__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14068_ net1239 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12170__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ team_02_WB.instance_to_wrap.top.pc\[31\] _06130_ vssd1 vssd1 vccd1 vccd1
+ _07539_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10334__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08560_ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] _04228_ _04226_ vssd1 vssd1
+ vccd1 vccd1 _04229_ sky130_fd_sc_hd__a21o_1
X_16709_ net1268 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
X_08491_ team_02_WB.instance_to_wrap.top.a1.data\[11\] net958 _04187_ vssd1 vssd1
+ vccd1 vccd1 _04188_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13036__C1 _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11062__A1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] net737 _04625_ _04627_
+ _04628_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_84_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09043_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] net884 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12345__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout309_A _06840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09558__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold421 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__A_N _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold454 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1120_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1218_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _04526_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
Xhold498 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\] net918 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ _05446_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout912 _04523_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout580_A _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 _04513_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_147_Left_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11117__A2 _06618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_2
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 _04500_ vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_2
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12080__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\] net761 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__a22o_1
Xfanout967 _02957_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_2
Xfanout978 _04281_ vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__buf_4
Xhold1110 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 _04431_ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09191__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1132 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ net1457 net1045 net992 team_02_WB.instance_to_wrap.ramaddr\[4\] vssd1 vssd1
+ vccd1 vccd1 _02598_ sky130_fd_sc_hd__a22o_1
XANTENNA__09730__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1143 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1165 team_02_WB.instance_to_wrap.ramload\[21\] vssd1 vssd1 vccd1 vccd1 net2527
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1187 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _04358_ _04360_ _04364_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__and3_1
Xhold1198 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07709_ _03302_ net425 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__xnor2_1
X_08689_ net1059 _04278_ _04315_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__or3_4
XANTENNA__13290__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ _06144_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_156_Left_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10548__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ net790 net551 _06166_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ _06097_ _06098_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__or2_1
X_13370_ net1057 team_02_WB.instance_to_wrap.top.ru.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _03014_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ net290 net2273 net567 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12255__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__A _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11457__A1_N net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net1235 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
XANTENNA__09549__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net269 net1978 net574 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11203_ net998 _06707_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__o21bai_1
X_12183_ net259 net2245 net576 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_165_Left_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11134_ net667 _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__or2_1
X_11065_ net398 _06448_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__nor2_1
X_15942_ clknet_leaf_6_wb_clk_i _02082_ _00750_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10016_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\] net684 _05528_ _05529_
+ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a2111oi_2
XANTENNA__09182__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09721__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15873_ clknet_leaf_102_wb_clk_i _02013_ _00681_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14824_ net1104 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ net1137 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_174_Left_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11967_ net340 net1922 net585 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
X_13706_ net1139 _03225_ _03226_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__nor3_1
XANTENNA__10095__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10918_ _06429_ _06431_ net401 vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__X _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14686_ net1127 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
X_11898_ net330 net2545 net486 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16425_ clknet_leaf_83_wb_clk_i _02560_ _01233_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dfrtp_1
X_13637_ net1562 net963 _03186_ _00018_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o211a_1
X_10849_ _04609_ net661 _06364_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a21o_2
XFILLER_0_144_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16356_ clknet_leaf_35_wb_clk_i _02496_ _01164_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09788__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13568_ team_02_WB.instance_to_wrap.top.lcd.nextState\[2\] net1052 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\]
+ _03103_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__and4b_1
XFILLER_0_82_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15307_ clknet_leaf_78_wb_clk_i team_02_WB.EN_VAL_REG _00120_ vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.testpc.en_latched sky130_fd_sc_hd__dfrtp_2
XANTENNA__15317__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12519_ net288 net1977 net447 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__mux2_1
X_16287_ clknet_leaf_61_wb_clk_i _02427_ _01095_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12165__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13499_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] _03063_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.lcd_en sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15238_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[29\]
+ _00051_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_183_Left_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15169_ net1145 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__09960__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ _03693_ net256 _03683_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a21o_1
X_09730_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] net923 net911 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a22o_1
XANTENNA__10307__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\] net728 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a221o_1
XANTENNA__09712__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08612_ net84 net1448 net957 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
X_09592_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\] net914 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08543_ net1547 net792 net651 _04188_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XANTENNA__13272__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout259_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08474_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nor2_2
XFILLER_0_119_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11035__A1 _05809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire609 _05270_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_2
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12075__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16242__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09026_ net944 _04505_ _04509_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__and3_4
XFILLER_0_143_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold240 team_02_WB.instance_to_wrap.top.a1.row2\[3\] vssd1 vssd1 vccd1 vccd1 net1602
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_X net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 team_02_WB.instance_to_wrap.ramaddr\[7\] vssd1 vssd1 vccd1 vccd1 net1613
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_02_WB.START_ADDR_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_02_WB.instance_to_wrap.ramaddr\[21\] vssd1 vssd1 vccd1 vccd1 net1635
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 team_02_WB.instance_to_wrap.ramaddr\[1\] vssd1 vssd1 vccd1 vccd1 net1646
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout720 _04384_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_8
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
Xfanout742 _04378_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_4
X_09928_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__inv_2
Xfanout753 net756 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_8
Xfanout764 _04373_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09164__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 _04369_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
Xfanout786 _04362_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09703__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09859_ net971 _05375_ net544 vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout797 net799 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
XFILLER_0_99_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12870_ _04423_ _07328_ _05877_ _05836_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_177_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ net300 net1821 net589 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10559__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ net1214 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
X_11752_ net286 net2440 net597 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10703_ _06219_ _06218_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__and2b_1
XANTENNA__10993__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__A_N net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14471_ net1182 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
X_11683_ _05970_ _07160_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_81_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13015__A2 _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16210_ clknet_leaf_77_wb_clk_i _02350_ _01018_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13422_ _03030_ _02765_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__nand2_1
XANTENNA_input91_A wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ team_02_WB.instance_to_wrap.top.pc\[25\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _06151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ clknet_leaf_48_wb_clk_i _02281_ _00949_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13353_ team_02_WB.instance_to_wrap.ramload\[15\] net1015 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[15\] sky130_fd_sc_hd__and2_1
X_10565_ net545 net387 _06081_ net391 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12304_ net359 net2266 net570 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ clknet_leaf_24_wb_clk_i _02212_ _00880_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13284_ net1633 net982 net964 _02991_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__a22o_1
X_10496_ _05380_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15023_ net1261 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
X_12235_ net2126 net331 net612 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
XANTENNA__10001__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ net323 net1884 net462 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ net948 _06618_ _06625_ net607 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__o211a_4
X_12097_ net1896 net318 net580 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15925_ clknet_leaf_31_wb_clk_i _02065_ _00733_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11048_ team_02_WB.instance_to_wrap.top.pc\[24\] _06267_ team_02_WB.instance_to_wrap.top.pc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__a21oi_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
XFILLER_0_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ clknet_leaf_30_wb_clk_i _01996_ _00664_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14807_ net1186 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10469__A _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15787_ clknet_leaf_15_wb_clk_i _01927_ _00595_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12999_ team_02_WB.instance_to_wrap.top.pc\[17\] _06192_ _07518_ vssd1 vssd1 vccd1
+ vccd1 _07519_ sky130_fd_sc_hd__a21boi_2
XANTENNA__10068__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14738_ net1185 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11999__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14669_ net1128 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16408_ clknet_leaf_100_wb_clk_i _02543_ _01216_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_08190_ _03906_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08969__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ clknet_leaf_47_wb_clk_i _02479_ _01147_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_191_Left_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10240__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12623__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09394__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13190__B2 _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07974_ _03601_ _03645_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__or3b_1
XANTENNA__09146__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ _05216_ _05217_ _05223_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nor4_2
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12859__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09644_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] net895 net891 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09575_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\] net773 net681 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\]
+ _05091_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _04213_ net1609 net849 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
XANTENNA__10059__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11195__A2_N net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08457_ _04158_ _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout710_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout808_A _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11702__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__and2b_1
XFILLER_0_190_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_154_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1240_X net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] net737 _05865_ _05866_
+ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10231__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _04295_ net945 _04505_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__and3_4
XFILLER_0_103_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10281_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\] net910 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10842__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09385__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ net278 net1810 net474 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__A2 _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09137__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 net551 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout561 net563 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_8
Xfanout572 net575 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_8
Xfanout583 _07209_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_4
X_13971_ net1252 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XFILLER_0_189_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout594 _07192_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_8
X_15710_ clknet_leaf_1_wb_clk_i _01850_ _00518_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11495__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _04489_ _06244_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__xnor2_1
X_16690_ clknet_leaf_70_wb_clk_i _02807_ _01414_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11495__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08685__C team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ clknet_leaf_124_wb_clk_i _01781_ _00449_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12853_ _05231_ _06194_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_202_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14984__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11247__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__or3b_2
XFILLER_0_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15572_ clknet_leaf_114_wb_clk_i _01712_ _00380_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12784_ _06918_ _06946_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14523_ net1077 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
X_11735_ net351 net1841 net600 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input94_X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14454_ net1109 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11666_ net511 _05511_ _06011_ _07151_ _05469_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13405_ _03300_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10617_ net551 _06133_ _06126_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__a21oi_4
X_14385_ net1221 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11597_ team_02_WB.instance_to_wrap.top.pc\[3\] net974 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\]
+ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16124_ clknet_leaf_20_wb_clk_i _02264_ _00932_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07623__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13336_ team_02_WB.instance_to_wrap.Wen _03297_ team_02_WB.instance_to_wrap.wb.curr_state\[0\]
+ _03301_ net2315 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a32o_1
X_10548_ _05231_ net406 vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16055_ clknet_leaf_120_wb_clk_i _02195_ _00863_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13267_ net1461 net983 net965 _02982_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a22o_1
XANTENNA__12443__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10479_ _05878_ _05880_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_94_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10752__A team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09376__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15006_ net1156 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
X_12218_ net1744 net262 net615 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__mux2_1
XANTENNA__09915__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _02953_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_write_i
+ sky130_fd_sc_hd__inv_2
XANTENNA__11059__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net248 net1701 net463 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XANTENNA__09128__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ clknet_leaf_36_wb_clk_i _02048_ _00716_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_07690_ _03385_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_108_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire609_A _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15839_ clknet_leaf_60_wb_clk_i _01979_ _00647_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\] net844 _04871_ _04873_
+ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_121_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08311_ _03997_ _03999_ _04018_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\] net826 net822 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12618__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08242_ _03949_ _03957_ _03941_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13222__A2_N net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08173_ _03849_ _03858_ _03891_ _03846_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11410__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12861__B _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12353__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_30_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__clkbuf_4
XANTENNA__13163__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09906__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout493_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XANTENNA__12910__A1 _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _03661_ _03673_ _03679_ _03659_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout660_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _03609_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or2_1
X_09627_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\] net700 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] net887 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__a22o_1
X_08509_ net1048 _04199_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12528__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\] net762 net748 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11520_ net946 _07007_ _07012_ net604 vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__o211a_4
XFILLER_0_136_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ net654 _06942_ _06946_ net665 _06945_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_152_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ net506 _05603_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__nand2_1
XANTENNA__10204__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ net1087 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
X_11382_ _05378_ _05931_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09070__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ net1026 _02891_ net1023 team_02_WB.instance_to_wrap.top.pc\[15\] vssd1 vssd1
+ vccd1 vccd1 _01496_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] net906 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_185_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10572__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12263__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input54_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _07358_ _07359_ _07434_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_76_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10264_ _05770_ _05776_ _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__nor3_1
XANTENNA__14979__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ net360 net2355 net479 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XANTENNA__12901__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10195_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\] net892 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\]
+ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_2
X_16742_ net1287 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
X_13954_ net1240 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XANTENNA__11468__B2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ _07366_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__or2_1
X_16673_ clknet_leaf_65_wb_clk_i _02790_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13209__A2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13885_ net1164 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15624_ clknet_leaf_16_wb_clk_i _01764_ _00432_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12836_ _04714_ _06143_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15555_ clknet_leaf_27_wb_clk_i _01695_ _00363_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12767_ _05558_ _05921_ _07282_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__or4_1
XANTENNA__12438__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14506_ net1178 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
X_11718_ net286 net1736 net601 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15486_ clknet_leaf_5_wb_clk_i _01626_ _00294_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12698_ net338 net1811 net431 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ net1173 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
X_11649_ net375 _06980_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or2_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09597__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput44 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
X_14368_ net1080 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
Xinput55 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09061__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput66 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
Xhold806 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xinput77 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ clknet_leaf_15_wb_clk_i _02247_ _00915_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold817 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13319_ _07183_ _02959_ team_02_WB.instance_to_wrap.top.pc\[0\] net1053 vssd1 vssd1
+ vccd1 vccd1 _03009_ sky130_fd_sc_hd__a2bb2o_1
Xinput88 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
Xhold828 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput99 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
Xhold839 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12173__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14299_ net1089 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
X_16038_ clknet_leaf_4_wb_clk_i _02178_ _00846_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11297__B _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ net165 net1043 net1035 net1451 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07811_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ _04419_ _04417_ net551 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07742_ _03431_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11459__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07673_ _03393_ _03394_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08875__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09412_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] net888 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09343_ _04853_ _04856_ _04858_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_36_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12348__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] net754 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a22o_1
X_08225_ _03905_ _03914_ _03927_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__and3_1
XFILLER_0_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1248_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ _03873_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10198__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12083__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10392__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ _03778_ _03780_ _03802_ _03806_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nand4_2
XFILLER_0_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout875_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09760__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net945 _04503_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__and3_4
XFILLER_0_199_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09512__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _06461_ _06462_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _03201_ _03202_ _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__or3_1
X_10882_ net416 _06388_ _06396_ net374 vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_211_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12621_ net1708 net292 net555 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10567__A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ clknet_leaf_84_wb_clk_i _00008_ _00153_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12552_ net290 net2194 net442 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XANTENNA__09291__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ _05918_ _05923_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15271_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[30\]
+ _00084_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12483_ net270 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] net559 vssd1
+ vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14222_ net1082 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11434_ net668 _06915_ _06927_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_151_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09043__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ net1216 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XANTENNA__16476__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11365_ net604 _06858_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_4_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_91_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13104_ _07466_ _07517_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13127__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10316_ _05829_ _05831_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_210_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14084_ net1091 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
X_11296_ net654 _06355_ _06797_ net419 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__o22ai_1
X_13035_ _07439_ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__xor2_1
X_10247_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] net767 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a22o_1
Xfanout1120 net1123 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_4
Xfanout1131 net1171 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__buf_2
XANTENNA__09751__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1142 net1146 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
X_10178_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net791 net650 _05694_
+ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a22oi_4
Xfanout1153 net1170 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_4
Xfanout1164 net1166 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_4
Xfanout1175 net1187 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_198_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1186 net1187 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_2
XANTENNA__08994__X _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14986_ net1142 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09503__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16725_ net1280 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13937_ net1233 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
XANTENNA__08857__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16656_ clknet_leaf_94_wb_clk_i _02775_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13868_ net1154 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15607_ clknet_leaf_115_wb_clk_i _01747_ _00415_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ _07340_ _07341_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__nor2_1
XANTENNA__12168__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13799_ net1426 _03284_ net961 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10477__A _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16587_ clknet_leaf_91_wb_clk_i _02706_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09050__B _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15538_ clknet_leaf_55_wb_clk_i _01678_ _00346_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09282__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15469_ clknet_leaf_48_wb_clk_i _01609_ _00277_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10764__X _06281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08010_ _03726_ _03727_ _03731_ _03719_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_71_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11800__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09034__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold647 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold658 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\] net702 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__a22o_1
XANTENNA__09990__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold669 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11129__B1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ net1047 _04200_ _04211_ net1009 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09892_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] net910 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a22o_1
XANTENNA__12631__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13207__A1_N _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ net152 net1042 net1034 net1422 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XANTENNA__16400__Q team_02_WB.instance_to_wrap.ramload\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04296_ _04302_ net932
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__and4_4
XFILLER_0_197_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07725_ _03413_ _03446_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__xor2_1
XANTENNA__08848__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12867__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A _07221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07656_ _03345_ _03361_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11490__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12078__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _03311_ _03312_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09326_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] net896 net943 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09273__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ _04764_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nor2_8
XANTENNA__12806__S _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11710__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08208_ _03897_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\] net746 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_78_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ _03849_ _03855_ _03857_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13109__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ net2385 net280 net639 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XANTENNA__09981__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__C team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10101_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\] net750 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__a22o_1
XANTENNA__12541__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _06172_ net652 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] net497
+ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ _05542_ _05544_ _05546_ _05548_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or4_1
X_14840_ net1197 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net1081 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XANTENNA__10849__X _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ net261 net2408 net480 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XANTENNA__08839__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ _03016_ net950 _03235_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__and3_1
X_16510_ clknet_leaf_27_wb_clk_i _02644_ _01317_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10934_ _06345_ _06447_ net371 vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16441_ clknet_leaf_43_wb_clk_i net1397 _01249_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_193_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ net1370 _04163_ net850 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
X_10865_ net368 _06041_ _06379_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12604_ net352 net1727 net438 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__mux2_1
X_16372_ clknet_leaf_14_wb_clk_i _02512_ _01180_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13584_ team_02_WB.instance_to_wrap.top.a1.row2\[16\] _03124_ _03129_ _03131_ _03138_
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a2111o_1
X_10796_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__inv_2
X_15323_ clknet_leaf_42_wb_clk_i _01466_ _00136_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ net358 net2500 net449 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
XANTENNA__11071__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11620__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15254_ clknet_4_6__leaf_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[13\]
+ _00067_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12466_ net331 net2193 net451 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205_ net1203 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ net1714 net314 net640 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15185_ net1140 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
X_12397_ net323 net2529 net458 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__mux2_1
XANTENNA__08989__X _04506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10031__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14136_ net1196 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
X_11348_ _06793_ _06847_ net370 vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__mux2_1
XANTENNA__12451__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ net1078 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
X_11279_ net668 _06768_ _06781_ net837 _06780_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__o221a_1
XANTENNA__09724__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _07446_ _07537_ _07444_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13193__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13284__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14969_ net1158 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
X_16708_ net1267 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_08490_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\] net979 vssd1 vssd1 vccd1
+ vccd1 _04187_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16639_ clknet_leaf_95_wb_clk_i _02758_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09255__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] net781 net741 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10935__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12626__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09042_ net944 _04528_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold411 team_02_WB.instance_to_wrap.top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 net1773
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10022__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold433 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold455 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16021__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\] net808 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\]
+ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__a221o_1
Xhold488 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net905 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12361__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout913 _04523_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_2
Xhold499 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1113_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 _04513_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09715__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout935 _02960_ vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
X_09875_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\] net749 net733 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__a22o_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 _04261_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
Xhold1100 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_4
XFILLER_0_209_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout573_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 _04177_ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_2
Xhold1111 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08826_ net133 net1040 net991 net1439 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
Xhold1133 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1166 team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net2528
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1177 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net846 _04360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout740_A _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] vssd1 vssd1 vccd1 vccd1
+ net2550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13275__B1 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1199 team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] vssd1 vssd1 vccd1 vccd1
+ net2561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout838_A _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07708_ _03400_ _03428_ _03429_ _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a22oi_4
X_08688_ net1060 _04315_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__or3b_1
XANTENNA__09494__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07639_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] _03335_ _03336_ _03361_ vssd1
+ vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _04494_ _06166_ _06126_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_76_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09246__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11589__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09309_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] net723 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__A2 _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _04886_ net406 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nor2_1
XANTENNA__12536__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11440__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12320_ net276 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\] net564 vssd1
+ vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10261__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ net261 net2324 net573 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__mux2_1
XANTENNA__10013__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11202_ _06184_ net653 net495 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] net497
+ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__a221o_1
XANTENNA__09954__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net248 net2305 net577 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__mux2_1
XANTENNA__11761__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__A _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net374 _06311_ _06342_ net379 _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__o221a_1
XANTENNA__10580__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15269__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11064_ net666 _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__nor2_1
X_15941_ clknet_leaf_28_wb_clk_i _02081_ _00749_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07592__C team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14987__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] net740 _05530_ _05531_
+ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a211o_1
X_15872_ clknet_leaf_17_wb_clk_i _02012_ _00680_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08985__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14823_ net1173 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13266__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11966_ net333 net2036 net584 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14754_ net1153 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
XANTENNA__09485__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10917_ net390 _06286_ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__a21oi_1
X_13705_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ _03222_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__and3_1
X_14685_ net1203 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
X_11897_ net337 net2035 net488 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13636_ _03023_ _03183_ _03185_ _03164_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__or4b_1
X_16424_ clknet_leaf_80_wb_clk_i _02559_ _01232_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10848_ net672 _06283_ _06284_ net670 _06363_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__a221o_1
XANTENNA__09237__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13567_ net1049 _03103_ _03104_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12446__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16355_ clknet_leaf_28_wb_clk_i _02495_ _01163_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10779_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__inv_2
X_15306_ clknet_leaf_69_wb_clk_i _01450_ _00119_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12518_ net277 net1904 net446 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__mux2_1
XANTENNA__10252__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16286_ clknet_leaf_5_wb_clk_i _02426_ _01094_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13498_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] _03019_ _03062_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12449_ net264 net2104 net452 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__mux2_1
X_15237_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[28\]
+ _00050_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_max_cap636_A _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10004__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09945__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15168_ net1145 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14119_ net1173 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XANTENNA__12181__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07990_ _03683_ _03693_ net256 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__nand3_2
X_15099_ net1080 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire541_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] net779 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ net85 net1513 net955 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_1
XANTENNA__08920__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09591_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\] net878 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08542_ team_02_WB.instance_to_wrap.top.a1.state\[2\] net793 vssd1 vssd1 vccd1 vccd1
+ _04224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08473_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ team_02_WB.instance_to_wrap.top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__or3b_1
XANTENNA__13025__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09228__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12864__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout321_A _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12356__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1063_A team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _04504_ _04516_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nor2_1
XANTENNA__10952__X _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1230_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09936__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net1592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13085__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold241 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net1603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 team_02_WB.instance_to_wrap.ramaddr\[14\] vssd1 vssd1 vccd1 vccd1 net1614
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 team_02_WB.instance_to_wrap.top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1 net1625
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12091__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09237__Y _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net712 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_8
Xfanout721 _04383_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_4
Xfanout732 _04381_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_8
X_09927_ net791 _05441_ _05443_ net650 vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a22oi_4
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout743 _04378_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 net756 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_8
Xfanout765 _04372_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 _04369_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
XANTENNA__16687__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ _05370_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_4
Xfanout787 _04362_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_8
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_4
X_08809_ net1510 net1041 net991 team_02_WB.instance_to_wrap.ramaddr\[22\] vssd1 vssd1
+ vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
X_09789_ _05298_ _05299_ _05301_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ net292 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\] net590 vssd1
+ vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XANTENNA__11259__C1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09467__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ net274 net2565 net598 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13650__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10702_ team_02_WB.instance_to_wrap.top.pc\[18\] _06188_ vssd1 vssd1 vccd1 vccd1
+ _06219_ sky130_fd_sc_hd__xnor2_1
X_14470_ net1212 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11682_ _04842_ _04861_ _05971_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__o211a_1
XANTENNA__09219__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ net1066 _03031_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10633_ _06128_ _06149_ _04490_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12266__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ clknet_leaf_126_wb_clk_i _02280_ _00948_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10234__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ net1533 net1016 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10564_ _04589_ net388 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__nor2_1
XANTENNA_input84_A wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12303_ net344 net2538 net571 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__mux2_1
X_16071_ clknet_leaf_40_wb_clk_i _02211_ _00879_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13283_ team_02_WB.instance_to_wrap.top.pc\[18\] net1053 _06759_ net935 vssd1 vssd1
+ vccd1 vccd1 _02991_ sky130_fd_sc_hd__a22o_1
X_10495_ _05993_ _06010_ _05992_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a21o_1
X_15022_ net1247 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
X_12234_ net1747 net334 net614 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
XANTENNA__07884__A team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12165_ net319 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\] net463 vssd1
+ vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net998 _06623_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13487__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12096_ net2343 net314 net582 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XANTENNA__13240__A_N _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15924_ clknet_leaf_4_wb_clk_i _02064_ _00732_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11047_ _06150_ net653 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] net496
+ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08902__B2 net2397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15855_ clknet_leaf_41_wb_clk_i _01995_ _00663_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14806_ net1084 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
X_15786_ clknet_leaf_39_wb_clk_i _01926_ _00594_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09458__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12998_ _07466_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__nand2b_1
X_14737_ net1229 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
X_11949_ net262 net1857 net587 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_157_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14668_ net1209 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16407_ clknet_leaf_105_wb_clk_i _02542_ _01215_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12176__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08418__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ team_02_WB.instance_to_wrap.top.a1.row1\[11\] _03110_ _03121_ team_02_WB.instance_to_wrap.top.a1.row1\[115\]
+ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14599_ net1182 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10225__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16338_ clknet_leaf_57_wb_clk_i _02478_ _01146_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09091__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16269_ clknet_leaf_49_wb_clk_i _02409_ _01077_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09918__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13190__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ _03647_ _03674_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__xnor2_2
X_09712_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] net676 _05213_ _05226_
+ _05228_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_126_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09697__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] net915 _05157_ _05159_
+ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a211o_1
XFILLER_0_184_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout271_A _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\] net749 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a22o_1
XANTENNA__09449__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net1048 _04211_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_26_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1180_A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ _04149_ _04150_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11008__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12086__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ _04094_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout703_A _04389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire429 _05623_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09082__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09621__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09008_ _04295_ net944 _04507_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10280_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] net894 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13469__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout551 _04356_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_4
Xfanout573 net574 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_8
X_13970_ net1252 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
Xfanout584 _07202_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_4
Xfanout595 _07192_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_4
XFILLER_0_189_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12921_ _07352_ _07440_ _07350_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11018__X _06530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15640_ clknet_leaf_122_wb_clk_i _01780_ _00448_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08685__D team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ _05231_ _06194_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_202_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11803_ net348 net2062 net593 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_14_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12783_ _06536_ _06569_ net416 vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__a21o_1
X_15571_ clknet_leaf_57_wb_clk_i _01711_ _00379_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14522_ net1089 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
X_11734_ net362 net2526 net600 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14453_ net1257 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
X_11665_ net511 _05511_ _05533_ _05556_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10207__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13404_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03016_
+ sky130_fd_sc_hd__nand3_1
X_10616_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] net996 _06127_ vssd1
+ vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__a21oi_1
X_14384_ net1226 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XANTENNA__09073__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input87_X net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11596_ net999 _07084_ net947 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09612__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16123_ clknet_leaf_30_wb_clk_i _02263_ _00931_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ _03296_ team_02_WB.instance_to_wrap.Ren team_02_WB.instance_to_wrap.wb.curr_state\[0\]
+ _03301_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _00014_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10547_ _05271_ net388 vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__nor2_1
XANTENNA__07623__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16054_ clknet_leaf_22_wb_clk_i _02194_ _00862_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13266_ net934 _02962_ _02981_ net1055 team_02_WB.instance_to_wrap.top.pc\[26\] vssd1
+ vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a32o_1
X_10478_ net547 net402 vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15005_ net1160 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
X_12217_ net1941 net267 net614 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__mux2_1
X_13197_ team_02_WB.instance_to_wrap.top.d_ready _03308_ _04286_ _04289_ vssd1 vssd1
+ vccd1 vccd1 _02953_ sky130_fd_sc_hd__or4_4
XANTENNA__08997__X _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12148_ net254 net1790 net465 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net1650 net238 net580 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XANTENNA__12132__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ clknet_leaf_27_wb_clk_i _02047_ _00715_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15838_ clknet_leaf_2_wb_clk_i _01978_ _00646_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15769_ clknet_leaf_123_wb_clk_i _01909_ _00577_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11803__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ _04009_ _04023_ _04017_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a21oi_2
X_09290_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] net928 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09851__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ net224 _03957_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12738__A2 _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _03806_ _03840_ _03847_ net227 _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a41o_1
XFILLER_0_12_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09603__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11598__X _07087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12634__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08811__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_99_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_28_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__clkbuf_4
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1026_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _03678_ _03657_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__and2b_1
XANTENNA__14150__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] net316 _03597_ vssd1 vssd1
+ vccd1 vccd1 _03610_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_50_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\] net787 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09557_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\] net920 _05072_ _05073_
+ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_65_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\] net979 vssd1 vssd1 vccd1
+ vccd1 _04200_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09488_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\] net843 _05002_ _05004_
+ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a211o_1
XFILLER_0_194_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09842__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08439_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04125_ vssd1 vssd1 vccd1
+ vccd1 _04144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ net416 _06504_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09055__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire226 _03936_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_1
X_10401_ _05648_ _05917_ _05647_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07605__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11381_ net795 _06874_ _06876_ net655 _06879_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__o221a_1
XANTENNA__12544__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10853__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13120_ _06834_ net232 _02890_ net976 _02888_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o221a_1
X_10332_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] net812 net808 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\]
+ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13051_ _07532_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__xnor2_1
X_10263_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\] net771 _05764_ _05778_
+ _05779_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_76_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12002_ net342 net2573 net480 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
X_10194_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\] net856 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__a22o_1
XANTENNA__08030__B2 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout370 net373 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout381 _06085_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_2
X_16741_ net1286 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
Xfanout392 _05856_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_2
X_13953_ net1238 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XANTENNA__13159__A_N net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ _05103_ _06188_ _07423_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__a21o_1
X_16672_ clknet_leaf_66_wb_clk_i _02789_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13884_ net1246 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15623_ clknet_leaf_40_wb_clk_i _01763_ _00431_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10587__X _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ _04672_ _06139_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15554_ clknet_leaf_117_wb_clk_i _01694_ _00362_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12766_ _05467_ _05514_ _05879_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__or4_1
XANTENNA__08097__B2 _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13090__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09833__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505_ net1216 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_11717_ net273 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\] net603 vssd1
+ vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12697_ net332 net2322 net430 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__mux2_1
X_15485_ clknet_leaf_13_wb_clk_i _01625_ _00293_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ net408 _07053_ _07132_ _07133_ net378 vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a221o_1
X_14436_ net1092 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XANTENNA__09046__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
XFILLER_0_126_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput45 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12454__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ net1115 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
X_11579_ net946 _07064_ _07068_ net604 vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__o211a_2
XANTENNA__14235__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput56 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_2
Xhold807 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
X_16106_ clknet_leaf_37_wb_clk_i _02246_ _00914_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput78 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
Xinput89 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
X_13318_ net1646 net982 net964 _03008_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__a22o_1
Xmax_cap526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold818 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ net1089 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
Xhold829 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_208_Right_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16037_ clknet_leaf_30_wb_clk_i _02177_ _00845_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13249_ team_02_WB.instance_to_wrap.top.pc\[31\] net1055 _06124_ _02968_ _02969_
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07810_ _03483_ _03529_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__xnor2_4
X_08790_ net1059 net648 _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a21o_1
X_07741_ _03461_ _03462_ _03436_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07672_ _03393_ _03394_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09411_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__clkinv_4
XANTENNA_wire507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12629__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\] net827 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\]
+ _04844_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_181_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09824__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] net743 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a22o_1
X_16699__1266 vssd1 vssd1 vccd1 vccd1 _16699__1266/HI net1266 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_16_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ net225 _03937_ _03939_ _03931_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a211o_1
XFILLER_0_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09037__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__Y _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08155_ _03827_ net227 _03820_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12364__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14145__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10198__A2 _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__inv_2
XANTENNA__10392__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16278__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11147__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout770_A _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__B2 _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\] net952 team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__and3b_2
XANTENNA__10370__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ _03601_ _03639_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ _06238_ _06463_ net974 vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_162_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10122__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09609_ net528 _05122_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10881_ _06394_ _06395_ net397 vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12539__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input101_A wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ net1754 net285 net552 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_195_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13072__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ net278 net1801 net442 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15212__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11502_ _05923_ _06005_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__xnor2_1
X_12482_ net263 net2516 net559 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
XANTENNA__09028__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15270_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[29\]
+ _00083_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11433_ net672 _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ net1122 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XANTENNA__12274__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14152_ net1104 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
X_11364_ _06197_ net652 _06837_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13103_ net1027 _02876_ net1025 team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1
+ vccd1 vccd1 _01499_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13127__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10315_ _05829_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_2
X_14083_ net1136 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11295_ _06579_ _06796_ net415 vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11138__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ _07353_ _07354_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__nand2_1
XANTENNA__08003__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10246_ net968 _05742_ _05761_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__o21a_1
XANTENNA__09200__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 net1119 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
Xfanout1121 net1123 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
XANTENNA__09155__Y _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1134 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_4
X_10177_ _05668_ _05693_ net551 vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__mux2_1
Xfanout1143 net1146 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_2
Xfanout1154 net1155 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
Xfanout1165 net1169 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_4
XANTENNA__13221__A2_N net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1176 net1179 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__buf_4
XANTENNA__12797__X _07321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1187 net1265 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_2
X_14985_ net1156 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
Xfanout1198 net1202 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16724_ net1279 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_105_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13936_ net1234 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10113__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ clknet_leaf_94_wb_clk_i _02774_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12449__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ net1163 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11206__X _06712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15606_ clknet_leaf_22_wb_clk_i _01746_ _00414_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12818_ _04172_ _04180_ _03317_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__a21oi_1
X_16586_ clknet_leaf_86_wb_clk_i _02705_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09267__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13798_ _03284_ _03285_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__nor2_1
XANTENNA__09806__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15537_ clknet_leaf_2_wb_clk_i _01677_ _00345_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12749_ _04906_ _04993_ _05038_ _05081_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15468_ clknet_leaf_126_wb_clk_i _01608_ _00276_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14419_ net1072 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16420__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12184__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ clknet_leaf_38_wb_clk_i _01539_ _00207_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold604 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold615 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold626 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_max_cap621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold659 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\] net762 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ net1541 _04437_ net930 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_09891_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\] net832 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08842_ net153 net1042 net1034 net1491 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_191_Right_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10352__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ _04359_ _04364_ _04370_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__and3_4
X_07724_ _03413_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10104__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _03363_ _03368_ _03376_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a21o_1
XANTENNA__12359__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout351_A _07126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1093_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09258__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13054__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07586_ team_02_WB.instance_to_wrap.top.pad.count\[0\] _03310_ vssd1 vssd1 vccd1
+ vccd1 _03312_ sky130_fd_sc_hd__or2_1
X_09325_ net533 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1260_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09256_ _04766_ _04768_ _04770_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__or4_4
XFILLER_0_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ _03911_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_43_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\] net763 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a22o_1
XANTENNA__12094__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1146_X net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _03849_ _03855_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09430__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _03788_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__or2_2
XANTENNA__14603__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] net770 net756 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a22o_1
XANTENNA__08023__D team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ team_02_WB.instance_to_wrap.top.pc\[24\] _06267_ vssd1 vssd1 vccd1 vccd1
+ _06590_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\] net835 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\]
+ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_164_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10343__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14770_ net1183 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
XANTENNA__09497__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ net266 net2618 net480 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XANTENNA__13293__B2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03235_
+ sky130_fd_sc_hd__a21o_1
X_10933_ net542 net387 _06316_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10578__A _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729__1357 vssd1 vssd1 vccd1 vccd1 net1357 _16729__1357/LO sky130_fd_sc_hd__conb_1
XFILLER_0_39_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12269__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16440_ clknet_leaf_45_wb_clk_i net1399 _01248_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
X_10864_ net367 _06047_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nand2_1
X_13652_ net1456 _04165_ net850 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XANTENNA__09249__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ net362 net2442 net438 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
X_16371_ clknet_leaf_56_wb_clk_i _02511_ _01179_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ _06303_ _06310_ net393 vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__mux2_1
X_13583_ _03132_ _03134_ _03137_ _03136_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or4b_1
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08990__B team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11901__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15322_ clknet_leaf_43_wb_clk_i _01465_ _00135_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07887__A team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12534_ net343 net2277 net447 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15253_ clknet_leaf_106_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[12\]
+ _00066_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12465_ net335 net2101 net452 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14204_ net1199 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11416_ net948 _06908_ _06913_ net607 vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__o211a_2
XANTENNA__09421__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12396_ net319 net2161 net458 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15184_ net1140 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14135_ net1209 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
X_11347_ _06308_ _06330_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__or2_1
XANTENNA__08775__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09607__A _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _05942_ _05980_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__xnor2_1
X_14066_ net1177 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
X_13017_ _07448_ _07536_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__or2_1
X_10229_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\] net855 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a22o_1
XANTENNA__10334__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 team_02_WB.instance_to_wrap.top.pad.button_control.debounce vssd1 vssd1 vccd1
+ vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_6_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14968_ net1198 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XANTENNA__11295__A0 _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16707_ net1349 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
X_13919_ net1228 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12179__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14899_ net1074 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16638_ clknet_leaf_95_wb_clk_i _02757_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13036__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16569_ clknet_leaf_87_wb_clk_i _02693_ _01376_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11811__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] net773 net761 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ _04626_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09660__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09041_ _04554_ _04555_ _04556_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or4_1
XFILLER_0_142_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10270__B2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09412__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold401 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold412 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12642__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold456 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold467 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] net914 net894 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout903 net905 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net917 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_8
Xfanout925 _04513_ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_4
XFILLER_0_0_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] net685 net681 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a22o_1
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_2
XANTENNA__10325__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout958 _04178_ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
Xhold1101 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 _04496_ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09191__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1123 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ net1446 net1041 net991 team_02_WB.instance_to_wrap.ramaddr\[6\] vssd1 vssd1
+ vccd1 vccd1 _02600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1134 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1167 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ net846 _04360_ _04364_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__and3_4
XANTENNA__13275__B2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1189 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07707_ _03364_ _03399_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__or2_1
XANTENNA__12089__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout733_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ net1059 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04316_ sky130_fd_sc_hd__nor2_1
XANTENNA__16466__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ _03356_ _03359_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] _03329_ vssd1
+ vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a2bb2o_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07569_ net1069 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout900_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1263_X net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11721__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10941__A1_N _04694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\] net691 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a22o_1
X_10580_ _04928_ net387 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\] net886 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12250_ net267 net2130 net573 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__mux2_1
XANTENNA__09403__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _06265_ _06706_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_170_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12181_ net254 net1876 net578 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__mux2_1
XANTENNA__12552__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _06296_ _06638_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold990 team_02_WB.instance_to_wrap.ramload\[4\] vssd1 vssd1 vccd1 vccd1 net2352
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15940_ clknet_leaf_35_wb_clk_i _02080_ _00748_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11063_ net416 _06569_ _06572_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__a21o_1
XANTENNA__11513__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] net772 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a22o_1
XANTENNA__11513__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09182__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ clknet_leaf_59_wb_clk_i _02011_ _00679_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12788__A _06508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14822_ net1205 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XANTENNA__13266__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13266__B2 team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ net1261 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
X_11965_ net335 net1972 net587 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] _03222_ net1636 vssd1
+ vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a21oi_1
X_10916_ net390 _06291_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14684_ net1201 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XANTENNA__09890__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net328 net2409 net489 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16423_ clknet_leaf_84_wb_clk_i _02558_ _01231_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] team_02_WB.instance_to_wrap.top.a1.row1\[101\]
+ _03184_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net667 _06344_ _06360_ net656 _06362_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16354_ clknet_leaf_117_wb_clk_i _02494_ _01162_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13206__A1_N _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ _03290_ _03115_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__and3_1
X_10778_ _06291_ _06293_ net368 vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__mux2_1
XANTENNA__09642__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15305_ clknet_leaf_67_wb_clk_i _01449_ _00118_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12517_ net283 net2365 net448 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16285_ clknet_leaf_13_wb_clk_i _02425_ _01093_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13497_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15236_ clknet_leaf_81_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[27\]
+ _00049_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12448_ net266 net1836 net453 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12970__B _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10771__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ net1145 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XANTENNA__12462__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ net255 net1697 net461 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14118_ net1213 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ net1074 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14049_ net1259 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10307__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11806__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ net86 net1433 _04261_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09590_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\] net825 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_50_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09072__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ _03291_ net792 _03319_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ team_02_WB.instance_to_wrap.top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_175_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload86_A clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12637__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09633__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16406__Q team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ _04519_ _04527_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1056_A team_02_WB.instance_to_wrap.top.ru.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12372__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__Y _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 team_02_WB.instance_to_wrap.top.a1.row2\[18\] vssd1 vssd1 vccd1 vccd1 net1593
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net1604 sky130_fd_sc_hd__dlygate4sd3_1
X_16728__1356 vssd1 vssd1 vccd1 vccd1 net1356 _16728__1356/LO sky130_fd_sc_hd__conb_1
Xhold253 team_02_WB.instance_to_wrap.ramaddr\[15\] vssd1 vssd1 vccd1 vccd1 net1615
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 team_02_WB.instance_to_wrap.ramaddr\[19\] vssd1 vssd1 vccd1 vccd1 net1626
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 team_02_WB.instance_to_wrap.top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1 net1637
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _04391_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
XANTENNA_fanout683_A _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 team_02_WB.instance_to_wrap.top.a1.row1\[113\] vssd1 vssd1 vccd1 vccd1 net1659
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
Xfanout722 _04383_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__clkbuf_4
X_09926_ _04417_ _05442_ net550 vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__mux2_1
Xfanout733 _04380_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_8
Xfanout744 _04378_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_2
Xfanout755 net756 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_4
XANTENNA__09164__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 _04372_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout777 _04367_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_4
X_09857_ _05359_ _05361_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__or3_1
Xfanout788 _04362_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 _04542_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_4
XANTENNA__11716__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ net1489 net1039 net993 team_02_WB.instance_to_wrap.ramaddr\[23\] vssd1 vssd1
+ vccd1 vccd1 _02617_ sky130_fd_sc_hd__a22o_1
X_09788_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\] net728 _05302_ _05304_
+ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__a211o_1
XANTENNA__15856__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ net932 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11750_ net288 net2002 net596 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__mux2_1
XANTENNA__09872__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ team_02_WB.instance_to_wrap.top.pc\[17\] _06190_ _06217_ vssd1 vssd1 vccd1
+ vccd1 _06218_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _05982_ _07165_ _07166_ _06019_ _04862_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__a311o_1
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ team_02_WB.instance_to_wrap.top.lcd.currentState\[2\] team_02_WB.instance_to_wrap.top.lcd.nextState\[2\]
+ net962 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10632_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net995 vssd1 vssd1 vccd1
+ vccd1 _06149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13351_ team_02_WB.instance_to_wrap.ramload\[13\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[13\] sky130_fd_sc_hd__and2_1
XFILLER_0_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10563_ _04631_ net403 vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__nor2_1
XANTENNA__15220__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ net340 net1827 net568 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16070_ clknet_leaf_7_wb_clk_i _02210_ _00878_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _05992_ _05993_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and2b_2
XANTENNA_input77_A wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13282_ net1626 net982 net964 _02990_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ net1168 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
XANTENNA__12282__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__B2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ net2512 net327 net614 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__mux2_1
X_12164_ net314 net1867 net464 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
XANTENNA__14998__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ net973 _06620_ _06621_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ net2103 net305 net583 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_207_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15923_ clknet_leaf_59_wb_clk_i _02063_ _00731_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11046_ _06151_ _06152_ _06233_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_207_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15854_ clknet_leaf_44_wb_clk_i _01994_ _00662_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10170__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14805_ net1200 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15785_ clknet_leaf_110_wb_clk_i _01925_ _00593_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12997_ _07467_ _07516_ _07469_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_203_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14736_ net1225 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ net265 net1825 net586 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_96_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11670__B1 _07150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12457__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14667_ net1125 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
X_11879_ net259 net2204 net486 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__mux2_1
X_16406_ clknet_leaf_100_wb_clk_i _02541_ _01214_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_184_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13618_ team_02_WB.instance_to_wrap.top.a1.row2\[11\] _03122_ _03124_ team_02_WB.instance_to_wrap.top.a1.row2\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a22o_1
XANTENNA__09615__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14598_ net1218 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10225__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16337_ clknet_leaf_1_wb_clk_i _02477_ _01145_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08969__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09091__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ net1051 _03290_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16268_ clknet_leaf_3_wb_clk_i _02408_ _01076_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13175__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15219_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[10\]
+ _00032_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12192__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ clknet_leaf_39_wb_clk_i _02339_ _01007_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07972_ _03684_ _03693_ _03680_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09146__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\] net722 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09642_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\] net872 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
XANTENNA__10161__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\] net785 net842 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout264_A _06595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\] net979 vssd1 vssd1 vccd1
+ vccd1 _04212_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13650__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09854__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _04149_ _04152_ _04150_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12367__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout431_A _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08386_ _04087_ _04089_ _04093_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout898_A _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09007_ _04313_ net944 _04507_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__and3_4
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09385__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09137__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\] net785 _05423_ _05425_
+ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__a211o_1
Xfanout552 net555 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_8
Xfanout563 _07219_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_8
Xfanout585 _07202_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
Xfanout596 _07191_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_8
X_12920_ _07353_ _07439_ _07354_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08896__B2 net2249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12851_ net520 _06192_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__15215__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13661__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ net352 net2597 net592 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_X clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15570_ clknet_leaf_54_wb_clk_i _01710_ _00378_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12782_ _07295_ _07302_ _07303_ _07305_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__and4_1
XANTENNA__09845__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14521_ net1090 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11733_ net357 net1921 net602 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XANTENNA__10586__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12277__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14058__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14452_ net1238 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
X_11664_ _05919_ _07146_ _07147_ _07149_ _07140_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__a41o_1
XFILLER_0_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ net2602 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1
+ vccd1 _03015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10615_ _03293_ _06130_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__xnor2_1
X_14383_ net1219 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11595_ team_02_WB.instance_to_wrap.top.pc\[3\] team_02_WB.instance_to_wrap.top.pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__xnor2_1
X_16122_ clknet_leaf_53_wb_clk_i _02262_ _00930_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13334_ _04243_ _04247_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__nand2_1
X_10546_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16053_ clknet_leaf_31_wb_clk_i _02193_ _00861_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13265_ _06523_ _02961_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__or2_1
X_10477_ _05440_ _05464_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15004_ net1147 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XANTENNA__09376__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ net1903 net258 net612 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16789__1333 vssd1 vssd1 vccd1 vccd1 _16789__1333/HI net1333 sky130_fd_sc_hd__conb_1
X_13196_ net1057 team_02_WB.instance_to_wrap.top.ru.state\[6\] team_02_WB.instance_to_wrap.Wen
+ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21o_4
XFILLER_0_209_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12147_ net238 net2097 net462 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09128__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ net1815 net246 net582 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
X_11029_ net416 _06536_ _06539_ net377 vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__a22o_1
X_15906_ clknet_leaf_116_wb_clk_i _02046_ _00714_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15837_ clknet_leaf_10_wb_clk_i _01977_ _00645_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15768_ clknet_leaf_123_wb_clk_i _01908_ _00576_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09836__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16727__1355 vssd1 vssd1 vccd1 vccd1 net1355 _16727__1355/LO sky130_fd_sc_hd__conb_1
XFILLER_0_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14719_ net1116 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XANTENNA__09300__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15699_ clknet_leaf_59_wb_clk_i _01839_ _00507_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_08240_ _03910_ _03942_ _03954_ _03955_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__or4_2
XFILLER_0_74_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08171_ _03778_ _03842_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__09367__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_11_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__clkbuf_4
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__12650__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1019_A _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ _03652_ _03655_ _03670_ _03672_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_182_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13320__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ net316 _03597_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1
+ vccd1 vccd1 _03609_ sky130_fd_sc_hd__a21oi_2
X_09625_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] net779 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a22o_1
X_09556_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] net916 net819 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\]
+ _05062_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09827__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08507_ team_02_WB.instance_to_wrap.top.a1.data\[7\] net958 vssd1 vssd1 vccd1 vccd1
+ _04199_ sky130_fd_sc_hd__or2_1
XFILLER_0_195_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12097__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] net742 net708 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\]
+ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout813_A _04521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ net1673 net1008 net981 _04143_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _04073_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10400_ _05912_ _05915_ _05691_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__o21ba_1
X_11380_ _06877_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10331_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\] net832 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09358__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ _07452_ _07453_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__and2b_1
X_10262_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\] net763 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12001_ net341 net2508 net481 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
X_10193_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\] net810 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\]
+ _05697_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__a221o_1
XANTENNA__12560__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
X_16740_ net1285 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_2
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_4
X_13952_ net1170 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
XFILLER_0_205_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10125__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15424__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ _07370_ _07422_ _07368_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09530__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16671_ clknet_leaf_66_wb_clk_i _02788_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13883_ net1253 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XFILLER_0_201_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11904__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15172__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15622_ clknet_leaf_9_wb_clk_i _01762_ _00430_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12834_ _04631_ _06134_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15553_ clknet_leaf_103_wb_clk_i _01693_ _00361_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12765_ _04567_ _06116_ _07283_ _07288_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14504_ net1105 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11716_ net290 net2013 net601 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
X_15484_ clknet_leaf_16_wb_clk_i _01624_ _00292_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12696_ net336 net2017 net433 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14435_ net1137 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
X_11647_ net390 _06285_ _07128_ net395 vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__o31a_1
XFILLER_0_142_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09597__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
X_14366_ net1189 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
Xinput35 gpio_in[20] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XFILLER_0_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput46 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
X_11578_ team_02_WB.instance_to_wrap.top.pc\[4\] net974 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\]
+ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__a221o_1
Xinput57 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ clknet_leaf_113_wb_clk_i _02245_ _00913_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput68 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold808 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16504__Q team_02_WB.START_ADDR_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13317_ team_02_WB.instance_to_wrap.top.pc\[1\] net1053 _07122_ net935 vssd1 vssd1
+ vccd1 vccd1 _03008_ sky130_fd_sc_hd__a22o_1
Xhold819 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ net504 net385 vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and2_1
Xinput79 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14297_ net1093 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
Xmax_cap538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_1
X_16036_ clknet_leaf_36_wb_clk_i _02176_ _00844_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13248_ _06124_ _02959_ _02966_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nor3_1
XFILLER_0_149_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12470__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10364__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _07048_ net232 _02937_ net976 _02939_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o221a_1
XFILLER_0_209_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09345__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__nand2_1
XANTENNA__10116__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _03356_ _03359_ _03388_ _03358_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_204_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11814__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _04915_ _04921_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__nor3_4
XFILLER_0_90_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09809__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09341_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\] net909 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\]
+ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_188_Left_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09272_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\] net787 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_115_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _03931_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12645__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ _03820_ _03827_ _03859_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__and3_1
XANTENNA__09588__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08424__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08085_ _03777_ _03804_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1136_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12380__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09760__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] _04502_ vssd1 vssd1
+ vccd1 vccd1 _04504_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout763_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10602__A1_N net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _03652_ _03655_ _03657_ _03659_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o211ai_1
XANTENNA__09512__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07869_ _03523_ _03562_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_162_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11724__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _05103_ _05122_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__or2_1
X_10880_ _06092_ _06096_ net373 vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\] net727 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_195_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13072__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16788__1332 vssd1 vssd1 vccd1 vccd1 _16788__1332/HI net1332 sky130_fd_sc_hd__conb_1
X_12550_ net280 net2184 net444 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11501_ net1660 net334 net639 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12555__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12481_ net266 net2159 net558 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__mux2_1
X_14220_ net1215 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
XANTENNA__12032__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _06011_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14151_ net1173 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
X_11363_ net975 _06209_ _06859_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__a31o_1
X_13102_ net978 _07423_ _02874_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__o31a_1
X_10314_ net395 net498 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14082_ net1191 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
X_11294_ net407 _06690_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_210_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15167__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ _07448_ _07536_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a21o_1
X_16726__1354 vssd1 vssd1 vccd1 vccd1 net1354 _16726__1354/LO sky130_fd_sc_hd__conb_1
XANTENNA__12290__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net969 _05742_ _05761_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10346__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1101 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
Xfanout1111 net1112 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_4
XANTENNA__10897__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] net648 _05692_ vssd1
+ vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a21o_1
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_2
XANTENNA__09751__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_201_Left_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1155 net1156 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
Xfanout1166 net1169 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_2
X_14984_ net1156 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
Xfanout1177 net1179 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1188 net1190 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
Xfanout1199 net1202 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_4
X_16723_ net1278 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_13935_ net1234 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
XANTENNA__09503__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16654_ clknet_leaf_94_wb_clk_i _02773_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13866_ net1162 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
XANTENNA__08509__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ clknet_leaf_40_wb_clk_i _01745_ _00413_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12817_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ team_02_WB.instance_to_wrap.top.a1.state\[0\] _03317_ vssd1 vssd1 vccd1 vccd1 _07340_
+ sky130_fd_sc_hd__and4b_1
X_16585_ clknet_leaf_86_wb_clk_i _02704_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13797_ net1641 _03282_ net961 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10110__Y _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15536_ clknet_leaf_30_wb_clk_i _01676_ _00344_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12748_ _04568_ _04609_ _04948_ _06113_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_210_Left_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12973__B _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10821__A1 _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12465__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15467_ clknet_leaf_14_wb_clk_i _01607_ _00275_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ net267 net2264 net432 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14418_ net1183 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15398_ clknet_leaf_8_wb_clk_i _01538_ _00206_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14349_ net1128 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold605 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold616 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold649 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16019_ clknet_leaf_58_wb_clk_i _02159_ _00827_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11809__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08910_ net1047 _04196_ _04208_ net1009 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a32o_1
X_09890_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\] net898 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ net154 net1043 net1035 net1453 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
XANTENNA__09742__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\] net685 net842 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a22o_1
X_07723_ _03416_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07654_ _03369_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09258__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07585_ net1859 _03311_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_A _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1086_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _04834_ _04836_ _04838_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__nor4_1
XFILLER_0_63_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09255_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] net922 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1253_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03858_ vssd1 vssd1 vccd1
+ vccd1 _03924_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12014__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_190_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09186_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] net751 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\]
+ _04697_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08769__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08137_ _03812_ _03850_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__xor2_2
XANTENNA__13995__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08068_ _03770_ _03787_ _03775_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__o21a_1
XANTENNA__09981__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout880_A _04538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11719__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_73_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] net901 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a22o_1
XANTENNA__09194__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_197_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ net257 net1543 net478 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _03015_ net950 _03234_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10932_ net417 _06438_ _06441_ net377 _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ net1595 _04167_ net850 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10863_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15223__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12602_ net356 net2396 net440 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16370_ clknet_leaf_54_wb_clk_i _02510_ _01178_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ team_02_WB.instance_to_wrap.top.a1.row1\[16\] _03111_ _03118_ team_02_WB.instance_to_wrap.top.a1.row2\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10794_ _06306_ _06309_ net368 vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15321_ clknet_leaf_45_wb_clk_i _01464_ _00134_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12533_ net339 net2021 net447 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
XANTENNA__12285__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15252_ clknet_leaf_104_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[11\]
+ _00065_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_191_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12464_ net326 net2400 net451 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__mux2_1
XANTENNA__15612__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14203_ net1075 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11415_ net994 _06910_ _06912_ _06837_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__a211o_1
X_15183_ net1140 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12395_ net314 net1531 net459 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08999__A team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10031__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14134_ net1121 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XANTENNA_input62_X net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ _05292_ net661 net658 _05293_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_120_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ net1229 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
X_11277_ _06037_ _06770_ _06778_ _06779_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__a211oi_1
X_13016_ _07449_ _07535_ _07450_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__o21a_1
XANTENNA__09724__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] net891 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 team_02_WB.instance_to_wrap.top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 net1364
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\] net911 net887 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11819__A0 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14967_ net1207 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
XANTENNA__10769__A _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13284__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16706_ net1348 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XANTENNA__10098__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13918_ net1167 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
X_14898_ net1183 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16637_ clknet_leaf_95_wb_clk_i _02756_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13849_ net1147 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13036__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11047__A1 _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16568_ clknet_leaf_90_wb_clk_i _02692_ _01375_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15519_ clknet_leaf_63_wb_clk_i _01659_ _00327_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12195__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16499_ clknet_leaf_127_wb_clk_i _02633_ _01306_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15292__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\] net834 net822 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\]
+ _04552_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_107_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold402 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10022__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09963__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold435 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold457 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11539__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09942_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\] net890 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold479 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout915 net917 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_8
X_16787__1331 vssd1 vssd1 vccd1 vccd1 _16787__1331/HI net1331 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_55_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout926 _04511_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_4
XANTENNA__09715__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout937 net938 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_1
X_09873_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\] net842 _05386_ _05387_
+ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_110_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout948 _04456_ vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_4
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout294_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 _04178_ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_2
Xhold1102 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ net1567 net1040 net991 team_02_WB.instance_to_wrap.ramaddr\[7\] vssd1 vssd1
+ vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1135 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net847 _04363_ _04368_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_116_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1157 team_02_WB.instance_to_wrap.top.pad.keyCode\[1\] vssd1 vssd1 vccd1 vccd1
+ net2519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1179 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _03399_ _03400_ net425 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a21boi_2
XANTENNA__10089__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ _04312_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or4_1
X_07637_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] _03329_ _03356_ _03359_ vssd1
+ vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_193_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout726_A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__A1 _05809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ team_02_WB.instance_to_wrap.top.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_192_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09100__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\] net755 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11589__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10261__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ net538 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\] net852 _04676_ _04685_
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ team_02_WB.instance_to_wrap.top.pc\[20\] _06264_ vssd1 vssd1 vccd1 vccd1
+ _06706_ sky130_fd_sc_hd__nor2_1
XANTENNA__10013__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12180_ net237 net1951 net576 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
XANTENNA__09954__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ net416 net412 vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nand2_1
Xhold980 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09706__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ net384 _06570_ _06571_ net377 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__a22o_1
XANTENNA__15218__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10013_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\] net728 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a22o_1
XANTENNA__09714__Y _05231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15870_ clknet_leaf_6_wb_clk_i _02010_ _00678_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_134_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1174 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XANTENNA__10589__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14752_ net1103 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ net327 net2542 net585 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
X_13703_ net2281 _03222_ _03224_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__o21a_1
X_10915_ net368 _06287_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14683_ net1084 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_11895_ net323 net2092 net486 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11912__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16422_ clknet_leaf_99_wb_clk_i _02557_ _01230_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_13634_ net1049 _03108_ _03135_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__o21ai_1
X_10846_ net381 net795 _06347_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__o31a_1
XFILLER_0_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16353_ clknet_leaf_104_wb_clk_i _02493_ _01161_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13565_ net1051 _03107_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_143_Left_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10777_ _05624_ net402 _06292_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08065__Y _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15304_ clknet_leaf_68_wb_clk_i _01448_ _00117_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12516_ net269 net1779 net449 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ clknet_leaf_16_wb_clk_i _02424_ _01092_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10252__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13496_ net191 net71 net104 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__and3b_1
XFILLER_0_136_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15235_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[26\]
+ _00048_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_140_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12447_ net260 net2295 net450 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__mux2_1
XANTENNA__11500__X _06994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__X _04694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09945__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15166_ net1144 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12378_ net236 net2269 net458 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14117_ net1113 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
X_11329_ net670 _06817_ _06829_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__a21bo_2
X_15097_ net1081 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
XANTENNA__09158__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14048_ net1080 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_152_Left_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15999_ clknet_leaf_62_wb_clk_i _02139_ _00807_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11268__A1 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _03313_ _04184_ net1577 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a21o_1
XANTENNA__09330__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _04169_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__or3b_1
XFILLER_0_82_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11822__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09023_ _04297_ _04500_ _04509_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12653__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout307_A _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__X _06908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09397__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold210 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13193__B2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 net169 vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 team_02_WB.START_ADDR_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16422__Q team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold243 net128 vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_02_WB.START_ADDR_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Left_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold265 team_02_WB.instance_to_wrap.ramaddr\[23\] vssd1 vssd1 vccd1 vccd1 net1627
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 team_02_WB.instance_to_wrap.top.a1.hexop\[1\] vssd1 vssd1 vccd1 vccd1 net1638
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout701 _04389_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_4
Xhold298 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 _04386_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
X_09925_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] _04330_ net649 team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a22o_1
Xfanout723 _04383_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_8
Xfanout734 _04380_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_4
Xfanout745 net748 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_8
Xfanout756 _04375_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_8
X_09856_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] net867 _05357_ _05372_
+ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a211o_1
Xfanout767 _04372_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_8
Xfanout778 _04367_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_4
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_4
X_08807_ net1549 net1040 net990 team_02_WB.instance_to_wrap.ramaddr\[24\] vssd1 vssd1
+ vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
X_09787_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] net780 net845 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout843_A _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08738_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04363_ _04365_ vssd1
+ vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__and3_4
XANTENNA__09321__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08669_ _04295_ _04296_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11732__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10700_ _06216_ _06215_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_159_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _04928_ _04947_ _04994_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ team_02_WB.instance_to_wrap.top.pc\[26\] _06147_ vssd1 vssd1 vccd1 vccd1
+ _06148_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ team_02_WB.instance_to_wrap.ramload\[12\] net1017 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[12\] sky130_fd_sc_hd__and2_1
XANTENNA__10234__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10562_ net542 net405 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13708__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12301_ net330 net2391 net568 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ _06731_ _02959_ team_02_WB.instance_to_wrap.top.pc\[19\] net1053 vssd1 vssd1
+ vccd1 vccd1 _02990_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12563__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ _05468_ _06009_ _05994_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09388__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15020_ net1165 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XANTENNA__13184__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ net1663 net324 net612 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__mux2_1
XANTENNA__11195__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ net306 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\] net465 vssd1
+ vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _06267_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ net2233 net298 net582 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__mux2_1
XANTENNA__13487__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ net672 _06533_ _06555_ net671 _06554_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__a221o_4
X_15922_ clknet_leaf_77_wb_clk_i _02062_ _00730_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_207_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11498__B2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15853_ clknet_leaf_49_wb_clk_i _01993_ _00661_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12447__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ net1153 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15784_ clknet_leaf_10_wb_clk_i _01924_ _00592_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12996_ team_02_WB.instance_to_wrap.top.pc\[15\] _06197_ _07515_ vssd1 vssd1 vccd1
+ vccd1 _07516_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09312__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14735_ net1220 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
X_11947_ net259 net1975 net584 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13423__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666_ net1176 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_11878_ net249 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] net487 vssd1
+ vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XANTENNA__08517__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16405_ clknet_leaf_100_wb_clk_i _02540_ _01213_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_13617_ _03164_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__nor2_1
X_16786__1330 vssd1 vssd1 vccd1 vccd1 _16786__1330/HI net1330 sky130_fd_sc_hd__conb_1
X_10829_ net545 net406 _06317_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a21o_1
X_14597_ net1175 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11422__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13548_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ _03289_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__and3_2
XFILLER_0_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16336_ clknet_leaf_23_wb_clk_i _02476_ _01144_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09091__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16267_ clknet_leaf_113_wb_clk_i _02407_ _01075_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10782__A _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13479_ team_02_WB.START_ADDR_VAL_REG\[19\] net1070 net1004 vssd1 vssd1 vccd1 vccd1
+ net202 sky130_fd_sc_hd__a21o_1
XANTENNA__12473__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09379__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15218_ clknet_leaf_104_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[9\]
+ _00031_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09918__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16198_ clknet_leaf_7_wb_clk_i _02338_ _01006_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07929__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15149_ net1144 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire644_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07971_ _03684_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11817__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] net766 net760 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__a22o_1
XANTENNA__11489__A1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] net907 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09572_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] net737 _05086_ _05088_
+ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a211o_1
XFILLER_0_210_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ team_02_WB.instance_to_wrap.top.a1.data\[3\] net958 vssd1 vssd1 vccd1 vccd1
+ _04211_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12648__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10957__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ _03307_ _04154_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10676__B _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_186_Right_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08385_ _04072_ _04077_ _04083_ _04078_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o31a_1
XFILLER_0_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout424_A _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1166_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10216__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09082__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12383__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11140__X _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ _04295_ _04501_ _04505_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__and3_4
XANTENNA__09909__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12913__A1 _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09790__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15823__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11727__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\] net721 net713 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__a221o_1
XANTENNA__12677__A0 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_6
Xfanout564 net567 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_8
Xfanout575 _07216_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_4
XANTENNA__13205__A1_N _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 _07202_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_8
Xfanout597 _07191_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_4
X_09839_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__inv_2
XANTENNA__10152__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12919__A2_N _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ net527 _06190_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11801_ net365 net2259 net592 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_202_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _06637_ _06696_ _06751_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__and4_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12558__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11101__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13243__A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14520_ net1196 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
X_11732_ net359 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] net602 vssd1
+ vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10586__B _06102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14451_ net1079 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
X_11663_ _07141_ _07148_ _05913_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15231__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13402_ net1623 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[31\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10207__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10614_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__inv_2
X_14382_ net1083 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
X_11594_ net794 _07074_ _07082_ net654 _07081_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__o221ai_4
XANTENNA__09073__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16121_ clknet_leaf_125_wb_clk_i _02261_ _00929_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13333_ net1057 net1661 net1053 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a21o_1
XANTENNA__11698__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ _05314_ net406 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12293__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ clknet_leaf_114_wb_clk_i _02192_ _00860_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13157__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ net1472 net983 net965 _02980_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__a22o_1
X_10476_ _05419_ net517 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15003_ net1133 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
XANTENNA__12904__A1 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12215_ net1704 net248 net614 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__mux2_1
X_13195_ net1027 _02952_ net1024 team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1
+ vccd1 vccd1 _01483_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_209_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09781__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net244 net2252 net464 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XANTENNA__09174__Y _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ net1656 net241 net582 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09533__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ _06385_ _06394_ net394 vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__mux2_1
X_15905_ clknet_leaf_103_wb_clk_i _02045_ _00713_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ clknet_leaf_17_wb_clk_i _01976_ _00644_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15767_ clknet_leaf_115_wb_clk_i _01907_ _00575_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12468__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ _07495_ _07498_ _07493_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14718_ net1190 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13066__A2_N net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15698_ clknet_leaf_18_wb_clk_i _01838_ _00506_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ net1091 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08170_ _03854_ _03860_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_172_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09064__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16319_ clknet_leaf_62_wb_clk_i _02459_ _01127_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_88_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__clkbuf_4
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08575__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
X_07954_ _03660_ _03664_ _03673_ _03676_ _03643_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_182_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07885_ _03576_ _03577_ _03598_ _03606_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _05129_ _05133_ _05137_ _05140_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] net900 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12378__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08506_ net2318 _04186_ _03319_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09486_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\] net784 net676 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ _04135_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1071_X net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout806_A _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ _04060_ _04070_ _04063_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09055__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08299_ _03983_ _04011_ _04013_ _03987_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_33_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10070__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10330_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\] _04529_ _04530_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a221o_1
XANTENNA__13139__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\] net787 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\]
+ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12000_ net330 net1839 net481 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09763__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\] net881 _05696_ _05708_
+ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_167_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout350 _07126_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_204_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 _07069_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09515__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13311__B2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_2
X_13951_ net1153 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
Xfanout394 net401 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_2
XANTENNA__15226__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _07369_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nand2_1
X_16670_ clknet_leaf_66_wb_clk_i _02787_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13882_ net1253 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ clknet_leaf_28_wb_clk_i _01761_ _00429_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12833_ _04631_ _06134_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12288__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15719__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11045__X _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12764_ _07284_ _07285_ _07286_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15552_ clknet_leaf_109_wb_clk_i _01692_ _00360_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09294__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ net278 net2015 net600 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
X_14503_ net1173 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15483_ clknet_leaf_34_wb_clk_i _01623_ _00291_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ net326 net2491 net431 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11920__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11646_ net389 _07089_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__nand2_1
X_14434_ net1191 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XANTENNA__09046__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1203 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_1
XFILLER_0_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput36 gpio_in[21] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_11577_ net1000 _07066_ net946 vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__o21ai_1
Xinput47 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput58 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16104_ clknet_leaf_24_wb_clk_i _02244_ _00912_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13316_ net1628 net984 net966 _03007_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__a22o_1
X_10528_ net501 net402 vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__and2_1
Xinput69 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
Xhold809 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ net1195 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
Xmax_cap528 net529 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16035_ clknet_leaf_9_wb_clk_i _02175_ _00843_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13247_ _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__inv_2
X_10459_ _04996_ _05041_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13178_ net229 _07501_ _02938_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__nand3_1
X_12129_ net307 net1873 net467 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XANTENNA__09506__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__B2 _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07670_ _03378_ _03387_ _03390_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__a211o_4
XFILLER_0_205_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15819_ clknet_leaf_15_wb_clk_i _01959_ _00627_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12198__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13605__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09340_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] net921 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_X clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\] net782 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11830__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08222_ _03921_ _03927_ _03901_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09037__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _03828_ _03858_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10052__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _03804_ _03777_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12661__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1129_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout491_A _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] _04502_ vssd1 vssd1
+ vccd1 vccd1 _04503_ sky130_fd_sc_hd__nor2_2
XFILLER_0_139_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ _03652_ _03655_ _03657_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o211a_1
X_16765__1309 vssd1 vssd1 vccd1 vccd1 _16765__1309/HI net1309 sky130_fd_sc_hd__conb_1
X_07868_ _03558_ _03565_ _03567_ _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_162_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ _05103_ _05122_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ _03490_ _03491_ net366 _03492_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout923_A _04513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09538_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\] net740 _05043_ _05047_
+ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09276__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\] net808 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\]
+ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11740__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ net946 _06989_ _06993_ net604 vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__o211a_2
X_12480_ net259 net2300 net556 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09028__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__Y _07221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11431_ _05465_ _05927_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13240__B _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10043__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14150_ net1213 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XANTENNA__08787__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ net1000 _06861_ _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1
+ vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__a2bb2o_1
X_13101_ net231 _02873_ _06761_ net234 vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ net408 net498 vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__nand2_1
X_14081_ net1259 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XANTENNA__12571__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ net407 _06794_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09736__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ net230 _07537_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08988__C team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net972 _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__or2_1
XANTENNA__09200__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16744__1289 vssd1 vssd1 vccd1 vccd1 _16744__1289/HI net1289 sky130_fd_sc_hd__conb_1
Xfanout1101 net1171 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1112 net1119 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_2
XANTENNA__10897__A2 _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] net997 _04329_ net1058
+ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a22o_1
Xfanout1123 net1131 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_2
XFILLER_0_206_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 net1146 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_4
Xfanout1156 net1170 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_4
XFILLER_0_206_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1167 net1169 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_4
X_14983_ net1142 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
XANTENNA__13296__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15541__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_2
XANTENNA__11915__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_4
X_16722_ net1277 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13934_ net1248 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08711__B2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16653_ clknet_leaf_95_wb_clk_i _02772_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13865_ net1162 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_202_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13599__A1 team_02_WB.instance_to_wrap.top.a1.row1\[58\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15604_ clknet_leaf_14_wb_clk_i _01744_ _00412_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12816_ team_02_WB.instance_to_wrap.top.edg2.flip1 _03299_ _04305_ vssd1 vssd1 vccd1
+ vccd1 _07339_ sky130_fd_sc_hd__a21oi_1
X_16584_ clknet_leaf_86_wb_clk_i _02703_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13796_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ _03280_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09267__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ clknet_leaf_44_wb_clk_i _01675_ _00343_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _07093_ _07094_ _07270_ _07074_ _07059_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_139_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10282__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15466_ clknet_leaf_37_wb_clk_i _01606_ _00274_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10821__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12678_ net258 net1905 net430 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08525__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14417_ net1226 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
X_11629_ net836 _07113_ _07115_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15397_ clknet_leaf_28_wb_clk_i _01537_ _00205_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10034__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09975__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ net1209 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold606 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold617 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold628 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ net1180 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XANTENNA__12481__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09727__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ clknet_leaf_55_wb_clk_i _02158_ _00826_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_08840_ net1479 net1044 net1036 net1441 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08771_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04296_ _04302_ net931
+ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__and4b_4
XFILLER_0_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11825__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _03410_ _03415_ net425 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__and3_1
XANTENNA_wire512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07653_ _03370_ _03371_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__or4_1
X_07584_ team_02_WB.instance_to_wrap.top.pad.count\[0\] _03310_ vssd1 vssd1 vccd1
+ vccd1 _03311_ sky130_fd_sc_hd__nand2_1
XANTENNA__09258__A2 _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09323_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\] net788 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a221o_1
XFILLER_0_192_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12656__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout337_A _06994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10273__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1079_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] net874 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08205_ _03862_ _03896_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] net710 _04699_ _04700_
+ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_190_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10025__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08136_ _03849_ _03855_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__and2_1
XANTENNA__09966__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A2 _04946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12391__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _03770_ _03775_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nor3_1
XANTENNA__14172__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_X clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1201_X net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14900__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13278__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\] net767 net679 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11735__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ net248 net2371 net480 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09497__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _06442_ _06443_ _06444_ net399 net382 vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__o221a_1
XFILLER_0_196_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ net390 _06043_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__or2_1
X_13650_ net1369 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] net851 vssd1 vssd1
+ vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
XANTENNA__09249__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ net359 net2418 net440 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
X_13581_ _03135_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03105_ vssd1
+ vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or3b_1
X_10793_ _06307_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12566__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13251__A _06365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15320_ clknet_leaf_42_wb_clk_i _01463_ _00133_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ net332 net2261 net446 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ net321 net2506 net450 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__mux2_1
X_15251_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[10\]
+ _00064_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10086__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14202_ net1090 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
X_11414_ net998 _06911_ _06833_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1
+ vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__a2bb2o_1
X_15182_ net1140 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
X_12394_ net305 net1995 net460 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14133_ net1241 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XANTENNA__08999__B team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ net422 _06313_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__nand2_1
XANTENNA__15178__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14064_ net1234 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XANTENNA_input55_X net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ net421 _06776_ _06358_ net655 vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_120_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13015_ team_02_WB.instance_to_wrap.top.pc\[27\] _06147_ _07534_ vssd1 vssd1 vccd1
+ vccd1 _07535_ sky130_fd_sc_hd__a21oi_1
X_10227_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] net912 net887 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a22o_1
XANTENNA__08932__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10158_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] net817 _04529_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ _05674_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a221o_1
XANTENNA__13269__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\] vssd1 vssd1 vccd1 vccd1
+ net1365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14966_ net1109 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
X_10089_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\] net774 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a22o_1
XANTENNA__09488__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16705_ net1347 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13917_ net1244 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
X_14897_ net1228 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16636_ clknet_leaf_95_wb_clk_i _02755_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13848_ net1148 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11047__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__A _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ clknet_leaf_87_wb_clk_i _02691_ _01374_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_13779_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] _03271_
+ net961 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_186_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10255__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15437__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15518_ clknet_leaf_5_wb_clk_i _01658_ _00326_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16498_ clknet_leaf_8_wb_clk_i _02632_ _01305_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09660__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15449_ clknet_leaf_125_wb_clk_i _01589_ _00257_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16764__1308 vssd1 vssd1 vccd1 vccd1 _16764__1308/HI net1308 sky130_fd_sc_hd__conb_1
XANTENNA__07713__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09412__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold425 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold436 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold447 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\] net828 _05447_ _05457_
+ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a211o_1
Xhold469 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout905 _04525_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__buf_4
XFILLER_0_110_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout916 net917 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_4
Xfanout927 _04511_ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
X_09872_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\] net785 net701 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\]
+ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 _02955_ vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_4
Xhold1103 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ net136 net1040 net991 net1424 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout287_A _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1136 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net846 _04363_ _04365_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__and3_4
Xhold1158 team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1 net2520
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10679__B _05785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07705_ net425 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08685_ net1058 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _04314_
+ sky130_fd_sc_hd__or4_1
XANTENNA__11286__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13680__B1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_A _07221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07636_ _03357_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_192_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__inv_2
XANTENNA__12386__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16743__1288 vssd1 vssd1 vccd1 vccd1 _16743__1288/HI net1288 sky130_fd_sc_hd__conb_1
X_09306_ net534 _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout719_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13071__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] net717 _04747_ _04752_
+ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_161_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1249_X net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\] net822 net810 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09403__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout990_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08119_ _03829_ _03836_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\] net785 net713 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ net423 net411 vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__nor2_1
Xhold970 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _06435_ _06439_ net393 vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__mux2_1
Xhold992 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14630__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\] net711 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a22o_1
XANTENNA__08914__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08914__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14820_ net1091 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XANTENNA__13246__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ net1117 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
X_11963_ net323 net2340 net584 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
XANTENNA__15234__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13702_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] _03222_ net1139 vssd1
+ vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10914_ net671 _06427_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__nand2_1
X_11894_ net317 net2583 net486 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
X_14682_ net1097 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09890__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16421_ clknet_leaf_95_wb_clk_i _02556_ _01229_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10845_ _04610_ net658 net664 _04611_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__o2bb2a_1
X_13633_ team_02_WB.instance_to_wrap.top.a1.row1\[109\] _03160_ _03168_ _03181_ _03182_
+ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12296__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11053__X _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ clknet_leaf_17_wb_clk_i _02492_ _01160_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10776_ net504 net402 vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__nand2_1
XANTENNA__08075__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13564_ _03104_ _03109_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09642__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15303_ clknet_leaf_68_wb_clk_i _01447_ _00116_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12515_ net261 net2309 net449 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08850__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16283_ clknet_leaf_33_wb_clk_i _02423_ _01091_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold990_X net2352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ team_02_WB.instance_to_wrap.top.ru.state\[4\] net1474 net1057 vssd1 vssd1
+ vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_dready sky130_fd_sc_hd__o21ba_1
XFILLER_0_137_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[25\]
+ _00047_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12446_ net249 net1846 net453 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08602__A0 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12377_ net245 net1808 net460 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__mux2_1
X_15165_ net1159 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11328_ net837 _06828_ _06827_ _06826_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__o211a_1
X_14116_ net1099 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15096_ net1172 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14047_ net1115 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
X_11259_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] net495 _06762_ net1001 net497
+ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ clknet_leaf_4_wb_clk_i _02138_ _00806_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14949_ net1174 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
XFILLER_0_210_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08470_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 _04169_
+ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_141_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09881__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16619_ clknet_leaf_90_wb_clk_i _02738_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10228__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09633__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14715__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ _04313_ net944 _04505_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__and3_4
XFILLER_0_127_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold200 net184 vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 team_02_WB.instance_to_wrap.top.a1.row1\[120\] vssd1 vssd1 vccd1 vccd1 net1573
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold222 team_02_WB.instance_to_wrap.ramaddr\[4\] vssd1 vssd1 vccd1 vccd1 net1584
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\] vssd1 vssd1 vccd1 vccd1
+ net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold244 _02596_ vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] vssd1 vssd1
+ vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 team_02_WB.instance_to_wrap.ramaddr\[2\] vssd1 vssd1 vccd1 vccd1 net1628
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold277 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold288 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09815__Y _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout702 _04389_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_2
Xhold299 team_02_WB.instance_to_wrap.top.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 net1661
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] _04330_ net649 team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a22o_1
Xfanout713 _04385_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_8
Xfanout724 _04383_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1209_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 _04380_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_8
Xfanout746 net748 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 net760 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
X_09855_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\] net814 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\]
+ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a221o_1
Xfanout768 _04372_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout571_A _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 _04367_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
X_08806_ net1476 net1040 net990 team_02_WB.instance_to_wrap.ramaddr\[25\] vssd1 vssd1
+ vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
X_09786_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] net744 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a22o_1
X_08737_ _04358_ _04360_ _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__and3_1
XANTENNA__11259__A2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__and2_2
XANTENNA__09872__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07619_ _03332_ _03335_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_159_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _03309_ net1003 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nor2_4
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ _06128_ _06146_ _04490_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_81_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11416__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09085__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ _06074_ _06077_ net370 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14625__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12300_ net334 net2208 net570 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13280_ net1553 net982 net964 _02989_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a22o_1
X_10492_ net511 _05511_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09388__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ net2433 net318 net612 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12162_ net296 net1861 net464 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
XANTENNA__15229__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ team_02_WB.instance_to_wrap.top.pc\[23\] _06266_ vssd1 vssd1 vccd1 vccd1
+ _06622_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ net1763 net308 net581 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ _06027_ _06531_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09454__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15921_ clknet_leaf_128_wb_clk_i _02061_ _00729_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_207_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08899__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__A2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15852_ clknet_leaf_126_wb_clk_i _01992_ _00660_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15282__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10170__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16763__1307 vssd1 vssd1 vccd1 vccd1 _16763__1307/HI net1307 sky130_fd_sc_hd__conb_1
XFILLER_0_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14803_ net1078 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
X_15783_ clknet_leaf_40_wb_clk_i _01923_ _00591_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12995_ _07470_ _07514_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__nor2_1
XANTENNA__11923__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15191__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14734_ net1076 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
X_11946_ net250 net2129 net586 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ net1210 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
X_11877_ net252 net1992 net487 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
X_16404_ clknet_leaf_100_wb_clk_i _02539_ _01212_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ _03103_ _03165_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a21o_1
X_10828_ net377 _06342_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09076__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ net1092 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XANTENNA__09615__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16335_ clknet_leaf_41_wb_clk_i _02475_ _01143_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08823__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ _03038_ _03057_ _03058_ _03040_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_99_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10759_ net975 _06275_ _06274_ _06253_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16266_ clknet_leaf_39_wb_clk_i _02406_ _01074_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13478_ team_02_WB.START_ADDR_VAL_REG\[18\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net201 sky130_fd_sc_hd__a21o_1
XANTENNA__13281__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15217_ clknet_leaf_105_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[8\]
+ _00030_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] sky130_fd_sc_hd__dfrtp_4
X_12429_ net318 net2296 net454 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16197_ clknet_leaf_29_wb_clk_i _02337_ _01005_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ net1157 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XANTENNA__10933__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _03690_ _03691_ _03686_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a21bo_1
X_15079_ net1263 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16742__1287 vssd1 vssd1 vccd1 vccd1 _16742__1287/HI net1287 sky130_fd_sc_hd__conb_1
X_09640_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\] net884 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10161__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\] net761 net705 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\]
+ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11833__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ _04210_ net1625 net849 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09854__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07612__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08453_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11134__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08384_ _04077_ _04086_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12664__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08814__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ net945 _04503_ _04507_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__and3_2
XFILLER_0_170_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11177__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_203_Right_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_A _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09907_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\] net681 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a22o_1
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_6
Xfanout565 net566 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 _07214_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_8
Xfanout587 _07202_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_4
X_09838_ _05348_ _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nor2_4
Xfanout598 _07191_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_6
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\] net826 net912 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\]
+ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11743__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11800_ net356 net2456 net594 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_202_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _06965_ _06982_ _07002_ _07056_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__and4_1
XANTENNA__11101__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09845__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ net344 net1894 net602 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14450_ net1183 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XANTENNA__09058__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11662_ net417 net500 _05914_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ net2344 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[30\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ net551 _06128_ _06129_ _06126_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a31o_2
X_11593_ net418 _06719_ _06921_ net376 _07073_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a221o_2
XANTENNA__12574__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14381_ net1126 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16120_ clknet_leaf_121_wb_clk_i _02260_ _00928_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10544_ _05356_ net386 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nor2_1
XANTENNA_input82_A wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13332_ _00008_ team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] vssd1 vssd1 vccd1
+ vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[4\] sky130_fd_sc_hd__or2_1
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11698__B _07183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ clknet_leaf_57_wb_clk_i _02191_ _00859_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13157__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ net517 _05419_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_134_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13263_ _02963_ _02979_ team_02_WB.instance_to_wrap.top.pc\[27\] net1056 vssd1 vssd1
+ vccd1 vccd1 _02980_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11168__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15002_ net1133 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XANTENNA__15648__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12214_ net1649 net255 net614 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13194_ net977 _02950_ _02951_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__o21a_1
XANTENNA__11918__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12145_ net242 net1794 net464 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XANTENNA__14090__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12076_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04452_ _06277_ _06279_
+ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__and4_4
X_11027_ net396 _06390_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__nand2_1
X_15904_ clknet_leaf_109_wb_clk_i _02044_ _00712_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10143__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ clknet_leaf_31_wb_clk_i _01975_ _00643_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15766_ clknet_leaf_21_wb_clk_i _01906_ _00574_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12978_ team_02_WB.instance_to_wrap.top.pc\[2\] _05836_ _07497_ vssd1 vssd1 vccd1
+ vccd1 _07498_ sky130_fd_sc_hd__a21o_1
XFILLER_0_188_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09836__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14717_ net1186 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929_ net322 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net482 vssd1
+ vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15697_ clknet_leaf_128_wb_clk_i _01837_ _00505_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14648_ net1195 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12484__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14265__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ net1078 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10603__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16318_ clknet_leaf_5_wb_clk_i _02458_ _01126_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16249_ clknet_leaf_123_wb_clk_i _02389_ _01057_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12356__A0 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_140_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09221__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11828__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_10_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__08710__B _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _03601_ _03663_ _03674_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_182_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13320__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07884_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] _03543_ _03575_ vssd1 vssd1
+ vccd1 vccd1 _03607_ sky130_fd_sc_hd__or3_1
XANTENNA__10134__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] net774 _05138_ _05139_
+ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a211o_1
XANTENNA__12659__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11416__X _06914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13344__A net2249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ _05064_ _05066_ _05068_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__or4_1
XANTENNA__09288__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08505_ net1048 _04185_ _04197_ _04198_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a31o_1
X_09485_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\] net734 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08990__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ _04137_ _04140_ _04139_ _04130_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12394__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ _04053_ _04074_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__xor2_1
XFILLER_0_163_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout701_A _04389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13188__A2_N net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08298_ _03978_ _03985_ _04012_ _03962_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09460__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13139__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16762__1306 vssd1 vssd1 vccd1 vccd1 _16762__1306/HI net1306 sky130_fd_sc_hd__conb_1
XFILLER_0_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\] net782 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a22o_1
XANTENNA__09212__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__A1 _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\] net835 net831 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10373__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_2
Xfanout351 _07126_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_204_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13311__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout373 _05857_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_2
X_13950_ net1243 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
Xfanout384 _06084_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10125__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net401 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_4
X_12901_ _05187_ _06192_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12569__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ net1250 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ clknet_leaf_36_wb_clk_i _01760_ _00428_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13254__A _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ _07350_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__nor2_1
XANTENNA__09279__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10597__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15551_ clknet_leaf_63_wb_clk_i _01691_ _00359_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12763_ _04782_ _04864_ _04995_ _05040_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__or4_1
XFILLER_0_185_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12822__A1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ net1212 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XFILLER_0_204_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11714_ net281 net2041 net603 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15482_ clknet_leaf_50_wb_clk_i _01622_ _00290_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12694_ net323 net2603 net430 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__mux2_1
X_14433_ net1256 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
X_11645_ _05902_ net660 _06116_ _07128_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__o2bb2a_1
X_16741__1286 vssd1 vssd1 vccd1 vccd1 _16741__1286/HI net1286 sky130_fd_sc_hd__conb_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ net1200 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09451__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_1
X_11576_ _06254_ _07065_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
X_16103_ clknet_leaf_38_wb_clk_i _02243_ _00911_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput48 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput59 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_13315_ team_02_WB.instance_to_wrap.top.pc\[2\] net1055 _07104_ net933 vssd1 vssd1
+ vccd1 vccd1 _03007_ sky130_fd_sc_hd__a22o_1
X_10527_ _06041_ _06043_ net389 vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14295_ net1208 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ clknet_leaf_117_wb_clk_i _02174_ _00842_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ _05127_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XANTENNA__09203__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246_ net934 _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13429__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ _07489_ _07490_ _07500_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__nand3b_1
X_10389_ _05832_ _05905_ _05829_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10364__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ net296 net2223 net468 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XANTENNA__13302__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ net303 net2438 net472 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux2_1
XANTENNA__10116__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12479__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15818_ clknet_leaf_32_wb_clk_i _01958_ _00626_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09809__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire502_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15749_ clknet_leaf_29_wb_clk_i _01889_ _00557_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\] net710 _04785_ _04786_
+ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a211o_1
XANTENNA__08493__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08221_ net226 _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08152_ _03828_ _03858_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__o31a_1
XANTENNA__13204__A1_N _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ _03771_ _03776_ _03787_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_184_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13219__A1_N net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10355__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] net952 vssd1 vssd1 vccd1
+ vccd1 _04502_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout484_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _03646_ _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nor2_1
XANTENNA__11304__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ _03558_ net329 _03565_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12389__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout749_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ net529 _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07798_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__inv_2
X_09537_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\] net845 _05048_ _05050_
+ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10985__X _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\] net922 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a22o_1
XANTENNA__15493__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10291__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ _04114_ _04121_ _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\] net718 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ net665 _06918_ _06925_ net654 _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ _06261_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13100_ _07368_ _07370_ _07422_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__and3_1
X_10312_ net395 net498 vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__or2_2
X_11292_ _06744_ _06793_ net370 vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__mux2_1
X_14080_ net1102 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10243_ _05754_ _05757_ _05758_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__or4_4
X_13031_ net1026 _02816_ net1024 team_02_WB.instance_to_wrap.top.pc\[30\] vssd1 vssd1
+ vccd1 vccd1 _01511_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10225__X _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10346__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_4
XANTENNA_input45_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ net504 _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__nor2_1
Xfanout1113 net1119 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_4
XFILLER_0_100_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15237__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1124 net1131 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_4
Xfanout1135 net1171 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_4
Xfanout1146 net1171 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09733__Y _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14982_ net1142 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
Xfanout1157 net1159 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_4
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_2
Xfanout1179 net1187 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_4
X_16721_ net1353 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_13933_ net1228 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XANTENNA__12299__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__A2 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16652_ clknet_leaf_94_wb_clk_i _02771_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ net1155 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13048__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15836__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15603_ clknet_leaf_56_wb_clk_i _01743_ _00411_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12815_ team_02_WB.instance_to_wrap.top.pc\[1\] team_02_WB.instance_to_wrap.top.testpc.en_latched
+ _07327_ _07336_ net1028 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a32o_1
XFILLER_0_186_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16583_ clknet_leaf_91_wb_clk_i _02702_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dfxtp_1
X_13795_ _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11931__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15534_ clknet_leaf_45_wb_clk_i _01674_ _00342_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12746_ _07269_ _07040_ _07023_ _07265_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__and4b_1
XANTENNA__09672__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07710__A team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15465_ clknet_leaf_107_wb_clk_i _01605_ _00273_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ net248 net2357 net432 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ net1226 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _05996_ net663 _06116_ _05878_ _07114_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__o221a_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15396_ clknet_leaf_36_wb_clk_i _01536_ _00204_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14347_ net1125 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11559_ team_02_WB.instance_to_wrap.top.pc\[5\] net974 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\]
+ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_133_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold607 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ net1213 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16017_ clknet_leaf_2_wb_clk_i _02157_ _00825_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13229_ net1576 net1021 net939 _05760_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11534__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11534__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08770_ _04302_ net847 _04364_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and3_4
XANTENNA__13287__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _03410_ net425 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07652_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nor2_1
XANTENNA__12002__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16761__1305 vssd1 vssd1 vccd1 vccd1 _16761__1305/HI net1305 sky130_fd_sc_hd__conb_1
XFILLER_0_192_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07583_ net2550 net1065 net34 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11841__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\] net728 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09253_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\] net808 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout232_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ _03917_ _03920_ _03903_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09184_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] net779 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ _04696_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a221o_1
XANTENNA__09415__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ _03852_ _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__and2b_1
XANTENNA__08769__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16141__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _03787_ _03321_ net1006 net1893 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13158__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1027_X net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout866_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\] net715 _04471_ _04484_
+ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a211o_1
X_16740__1285 vssd1 vssd1 vccd1 vccd1 _16740__1285/HI net1285 sky130_fd_sc_hd__conb_1
X_07919_ _03601_ _03639_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__and2b_1
X_08899_ net27 net1033 net989 net2572 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_197_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ _06323_ _06340_ net391 vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_104_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10861_ _06375_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__inv_2
XFILLER_0_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11751__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14628__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net342 net2280 net439 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ net1052 _03115_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__nand2_1
XANTENNA__09654__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10792_ _05271_ net404 vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ net334 net1973 net449 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15239__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15250_ clknet_leaf_106_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[9\]
+ _00063_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09406__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12462_ net317 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\] net450 vssd1
+ vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ net1099 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
X_11413_ team_02_WB.instance_to_wrap.top.pc\[12\] _06259_ vssd1 vssd1 vccd1 vccd1
+ _06911_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12582__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ net1140 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12393_ net296 net2108 net460 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14132_ net1239 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
X_11344_ _05935_ _06843_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09176__B _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14063_ net1224 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
X_11275_ _05980_ _06110_ _06775_ _06104_ _06777_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ _07451_ _07533_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__nor2_1
XANTENNA__09185__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] net895 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a22o_1
XANTENNA__11926__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] net927 net923 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a22o_1
Xhold4 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\] vssd1 vssd1
+ vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14965_ net1242 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
X_10088_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] net760 net732 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a22o_1
XANTENNA__11227__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16704_ net1346 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
X_13916_ net1252 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14896_ net1232 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
XANTENNA__09893__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16635_ clknet_leaf_95_wb_clk_i _02754_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13847_ net1138 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XANTENNA__14538__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16566_ clknet_leaf_89_wb_clk_i _02690_ _01373_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13778_ _03271_ _03272_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_44_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09645__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_X clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16526__Q net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15517_ clknet_leaf_13_wb_clk_i _01657_ _00325_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12729_ _06585_ _06792_ _06817_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__or4b_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16497_ clknet_leaf_127_wb_clk_i _02631_ _01304_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15448_ clknet_leaf_122_wb_clk_i _01588_ _00256_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12492__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15379_ clknet_leaf_83_wb_clk_i _01519_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold404 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold459 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09940_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\] net874 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a22o_1
XANTENNA__11507__B2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout906 _04524_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] net741 net721 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a22o_1
Xfanout917 _04518_ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 _04511_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_8
Xfanout939 _02954_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
XANTENNA__11836__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ net137 net1045 net992 net1378 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
Xhold1104 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 team_02_WB.instance_to_wrap.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net2477
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1137 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net847 _04368_ _04370_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__and3_4
Xhold1148 team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net2510
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ _03420_ _03425_ _03426_ _03393_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a22o_1
XANTENNA__10041__A _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_179_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09884__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] _03324_ _03328_ vssd1 vssd1
+ vccd1 vccd1 _03358_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12667__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout447_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__Y _04346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07566_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 _03306_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09636__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09305_ net970 _04821_ net543 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o21a_1
XANTENNA__09100__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10246__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09236_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] net765 net685 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08733__X _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09167_ _04678_ _04680_ _04682_ _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__or4_1
XANTENNA__13097__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ _03793_ _03830_ _03831_ _03790_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_2_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09098_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] net777 net729 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\]
+ _04612_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_170_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout983_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ _03763_ _03764_ _03769_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__a21o_1
Xhold960 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _06440_ _06444_ net394 vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__mux2_1
Xhold982 team_02_WB.instance_to_wrap.ramload\[30\] vssd1 vssd1 vccd1 vccd1 net2344
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _05516_ _05520_ _05524_ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10182__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16037__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14750_ net1189 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_11962_ net319 net2210 net584 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XANTENNA__09875__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _03222_ _03223_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__nor2_1
X_10913_ _04695_ _06031_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12577__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ net1097 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
X_11893_ net314 net2532 net487 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XANTENNA__11481__S net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16420_ clknet_leaf_80_wb_clk_i _02555_ _01228_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13632_ team_02_WB.instance_to_wrap.top.a1.row1\[13\] _03109_ _03114_ _03117_ team_02_WB.instance_to_wrap.top.a1.row1\[61\]
+ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__a32o_1
X_10844_ net424 _06354_ _06357_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09627__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16351_ clknet_leaf_59_wb_clk_i _02491_ _01159_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13563_ net1050 net1051 _03290_ _03103_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10775_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08075__B _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ clknet_leaf_68_wb_clk_i _01446_ _00115_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ net265 net2265 net448 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16282_ clknet_leaf_53_wb_clk_i _02422_ _01090_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13494_ team_02_WB.instance_to_wrap.top.d_ready _04286_ _04289_ team_02_WB.instance_to_wrap.top.ru.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_read_i sky130_fd_sc_hd__o31a_1
XFILLER_0_192_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15189__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15233_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[24\]
+ _00046_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ net255 net1734 net452 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15164_ net1144 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12376_ net241 net2311 net460 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__mux2_1
X_16760__1304 vssd1 vssd1 vccd1 vccd1 _16760__1304/HI net1304 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_97_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14115_ net1136 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
X_11327_ _05939_ _05988_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15095_ net1074 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ net1189 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
X_11258_ _06761_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\] net772 _05724_ _05725_
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a211o_1
XANTENNA__10173__A0 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net545 net398 _06692_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_128_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15997_ clknet_leaf_13_wb_clk_i _02137_ _00805_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14948_ net1093 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09866__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09330__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879_ net1109 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14268__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16618_ clknet_leaf_90_wb_clk_i _02737_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09618__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16549_ clknet_leaf_88_wb_clk_i _02673_ _01356_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13900__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_75_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ _04313_ net945 _04505_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and3_4
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09368__Y _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09397__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold201 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 net117 vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 team_02_WB.instance_to_wrap.top.a1.row1\[112\] vssd1 vssd1 vccd1 vccd1 net1596
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold245 net109 vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14731__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold256 team_02_WB.instance_to_wrap.ramstore\[20\] vssd1 vssd1 vccd1 vccd1 net1618
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 team_02_WB.instance_to_wrap.ramaddr\[17\] vssd1 vssd1 vccd1 vccd1 net1629
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 team_02_WB.instance_to_wrap.ramaddr\[6\] vssd1 vssd1 vccd1 vccd1 net1640
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net513 vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__inv_2
XANTENNA__09149__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold289 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout703 _04389_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout714 _04385_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 _04382_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_4
Xfanout736 _04380_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_4
X_09854_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] net911 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a22o_1
XANTENNA__10164__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout758 net760 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_8
Xfanout769 _04371_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_84_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08805_ net1402 net1045 net992 team_02_WB.instance_to_wrap.ramaddr\[26\] vssd1 vssd1
+ vccd1 vccd1 _02620_ sky130_fd_sc_hd__a22o_1
X_09785_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\] net783 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout564_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__and3b_2
XANTENNA__10977__Y _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09321__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] _03329_ _03338_ _03340_ vssd1
+ vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _04250_ _04251_ _04253_ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__or4_1
XFILLER_0_193_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07549_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1
+ _03290_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1261_X net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10560_ _06075_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or2_1
XANTENNA__13169__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\] net701 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10491_ net511 _05511_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_20_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09719__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09388__A2 _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net2290 net314 net614 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ net309 net2040 net463 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ _04494_ net653 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] net496
+ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__a221o_1
XANTENNA__09735__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net2206 net302 net583 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold790 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11329__X _06830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _06551_ _06552_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__or3b_1
X_15920_ clknet_leaf_23_wb_clk_i _02060_ _00728_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10155__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09560__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ clknet_leaf_14_wb_clk_i _01991_ _00659_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15245__Q team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14802_ net1184 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
X_15782_ clknet_leaf_6_wb_clk_i _01922_ _00590_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09848__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _07471_ _07513_ _07472_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09312__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ net1126 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
X_11945_ net252 net1644 net587 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12100__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14664_ net1111 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ net238 net2096 net486 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16403_ clknet_leaf_106_wb_clk_i _02538_ _01211_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__B1 _06901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13615_ team_02_WB.instance_to_wrap.top.lcd.nextState\[4\] _03105_ _03113_ _03165_
+ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a32o_1
X_10827_ net421 _06313_ _06329_ net379 vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14595_ net1136 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16334_ clknet_leaf_46_wb_clk_i _02474_ _01142_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13546_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _03061_ _03092_ net1068
+ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_99_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10758_ _06242_ _06246_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_99_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16265_ clknet_leaf_116_wb_clk_i _02405_ _01073_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13477_ team_02_WB.START_ADDR_VAL_REG\[17\] _04260_ vssd1 vssd1 vccd1 vccd1 net200
+ sky130_fd_sc_hd__and2_1
X_10689_ _03294_ _06203_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15216_ clknet_leaf_98_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[7\]
+ _00029_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09379__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ net312 net2472 net455 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__mux2_1
X_16196_ clknet_leaf_35_wb_clk_i _02336_ _01004_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ net1157 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
X_12359_ net308 net1852 net563 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15078_ net1246 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14029_ net1122 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XANTENNA__13167__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10146__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16352__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09570_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] net777 net713 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__a22o_1
X_08521_ _04171_ _04208_ _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08452_ _04145_ _04153_ _04148_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12010__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08383_ _04082_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__or2_1
XANTENNA__14726__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1054_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _04297_ _04500_ _04503_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__and3_2
XFILLER_0_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12680__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09790__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout681_A _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\] net761 net745 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__a22o_1
XANTENNA__11149__X _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10137__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 _04498_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_4
Xfanout555 _07227_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_4
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_6
XANTENNA__09542__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] net742 _05350_ _05352_
+ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__a2111o_1
Xfanout577 _07214_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_4
Xfanout588 net591 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_6
Xfanout599 _07191_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_4
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\] net864 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08719_ net1061 _04277_ _04323_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_202_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09699_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] net720 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11730_ net338 net2312 net601 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ _05624_ _05646_ _05920_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__or3b_1
XFILLER_0_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ net2510 net1011 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[29\]
+ sky130_fd_sc_hd__and2_1
X_10612_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net995 vssd1 vssd1 vccd1
+ vccd1 _06129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14380_ net1209 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11592_ net665 _07076_ _07078_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13331_ net1586 _03013_ _03010_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[3\]
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_181_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10543_ net390 _06055_ _06056_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16050_ clknet_leaf_76_wb_clk_i _02190_ _00858_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input75_A wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ _06490_ _02962_ _02959_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a21o_1
X_10474_ _05314_ _05334_ _05377_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11168__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15001_ net1148 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
X_12213_ net1737 net239 net613 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12590__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13193_ net230 _02949_ team_02_WB.instance_to_wrap.top.pc\[2\] net233 vssd1 vssd1
+ vccd1 vccd1 _02951_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10376__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ net643 _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nand2_4
XANTENNA__09781__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12075_ net346 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\] net470 vssd1
+ vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XANTENNA__10404__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15903_ clknet_leaf_61_wb_clk_i _02043_ _00711_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09533__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ net397 _06395_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__or2_1
XANTENNA__11934__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ clknet_leaf_50_wb_clk_i _01974_ _00642_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11628__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15765_ clknet_leaf_31_wb_clk_i _01905_ _00573_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12977_ _07334_ _07496_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__and2b_1
XANTENNA__11235__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11928_ net318 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\] net482 vssd1
+ vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__mux2_1
X_14716_ net1192 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
X_15696_ clknet_leaf_22_wb_clk_i _01836_ _00504_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14647_ net1186 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
X_11859_ net313 net2291 net491 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14578_ net1183 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XANTENNA__10603__A1 _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16317_ clknet_leaf_4_wb_clk_i _02457_ _01125_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13529_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _03061_ _03080_ _03089_
+ net1068 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16248_ clknet_leaf_114_wb_clk_i _02388_ _01056_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Left_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
X_16179_ clknet_leaf_52_wb_clk_i _02319_ _00987_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__10367__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12005__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _03663_ _03674_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nand2_1
XANTENNA__10119__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07883_ net316 _03597_ _03578_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11844__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] net770 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_158_Left_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09553_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\] net942 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\]
+ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A _06595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08504_ team_02_WB.instance_to_wrap.top.a1.row1\[16\] net849 vssd1 vssd1 vccd1 vccd1
+ _04198_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09484_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\] net698 net686 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ _04139_ _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__and2b_1
XFILLER_0_175_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12675__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1171_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13360__A net2520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ _04075_ _04076_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08297_ _03306_ _03746_ _03964_ _03972_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__or4_1
XANTENNA__15272__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] net929 net901 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09763__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout330 _07013_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_2
Xfanout341 _07030_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11858__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout352 _07126_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09515__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout363 _07107_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
XANTENNA__11754__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 net400 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_2
XANTENNA__08723__B1 _04346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ _07371_ _07419_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__and2_1
X_13880_ net1250 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _04589_ _06131_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15550_ clknet_leaf_5_wb_clk_i _01690_ _00358_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12762_ _05126_ _05210_ _05293_ _05379_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__or4_1
XFILLER_0_185_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ net1172 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ net271 net2257 net603 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XANTENNA__08067__C _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ clknet_leaf_125_wb_clk_i _01621_ _00289_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12693_ net319 net2422 net430 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__mux2_1
XANTENNA__12585__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08635__Y _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14432_ net1081 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11644_ _07129_ _04462_ _06114_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_5_0_wb_clk_i_X clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14363_ net1084 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ team_02_WB.instance_to_wrap.top.pc\[3\] team_02_WB.instance_to_wrap.top.pc\[2\]
+ team_02_WB.instance_to_wrap.top.pc\[4\] vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__a21oi_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XFILLER_0_91_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16102_ clknet_leaf_8_wb_clk_i _02242_ _00910_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput38 wb_rst_i vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_13314_ net1429 net983 net965 _03006_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10526_ _05995_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__or2_1
XANTENNA__10061__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput49 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
X_14294_ net1084 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11929__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16033_ clknet_leaf_101_wb_clk_i _02173_ _00841_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13245_ _06365_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
X_10457_ _05972_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__nor2_1
XANTENNA__10349__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__C1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13176_ _07398_ _07400_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__xnor2_1
X_10388_ _05878_ _05903_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08962__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ net308 net2591 net469 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09923__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ net295 net2473 net471 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__mux2_1
X_11009_ _06122_ _06517_ _06520_ _06509_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__a211o_1
X_15817_ clknet_leaf_110_wb_clk_i _01957_ _00625_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_16797_ net1341 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11077__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15748_ clknet_leaf_34_wb_clk_i _01888_ _00556_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12495__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ clknet_leaf_61_wb_clk_i _01819_ _00487_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14276__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ _03916_ _03926_ _03920_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_138_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ _03849_ _03855_ _03857_ _03826_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_151_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08082_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16690__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13339__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ net1058 net952 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ _03614_ _03637_ _03617_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_149_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout477_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07866_ _03558_ _03563_ _03564_ net329 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__nand4_1
X_09605_ net971 net628 net544 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_162_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07797_ _03491_ _03514_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__xnor2_2
X_09536_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\] net776 _05051_ _05052_
+ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a211o_1
XFILLER_0_168_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12265__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09130__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] net820 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\]
+ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10918__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14186__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_A _04524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ _04125_ _03321_ net1008 net1611 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_163_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09398_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\] net787 _04911_ _04912_
+ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_175_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08349_ _04047_ _04049_ _04058_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__or3_1
XFILLER_0_190_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10219__A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14914__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10043__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09984__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ team_02_WB.instance_to_wrap.top.pc\[14\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _06860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ _05811_ _05817_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__nor3_1
XANTENNA__11749__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ _05187_ net404 _06332_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_91_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13030_ net977 _02815_ _07547_ _07544_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__o211a_1
XANTENNA__09736__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\] net826 net900 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\]
+ _05745_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_210_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1103 net1110 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
X_10173_ _05671_ net622 net968 vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1114 net1119 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__buf_2
Xfanout1125 net1131 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_4
XFILLER_0_100_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1136 net1138 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_4
XANTENNA_input38_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1149 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__buf_4
XANTENNA__10889__A _05809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14981_ net1156 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
Xfanout1158 net1159 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_4
XANTENNA__13296__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_2
X_16720_ net1352 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XANTENNA__13265__A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13932_ net1233 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16651_ clknet_leaf_94_wb_clk_i _02770_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13863_ net1149 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
XANTENNA__08711__A3 _04339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12814_ team_02_WB.instance_to_wrap.top.testpc.en_latched team_02_WB.instance_to_wrap.top.i_ready
+ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__nand2_1
X_15602_ clknet_leaf_54_wb_clk_i _01742_ _00410_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13794_ net2122 _03280_ net961 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__o21ai_1
X_16582_ clknet_leaf_92_wb_clk_i _02701_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09121__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12745_ _06609_ _07267_ _07268_ _06643_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__or4b_1
X_15533_ clknet_leaf_47_wb_clk_i _01673_ _00341_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10282__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15464_ clknet_leaf_11_wb_clk_i _01604_ _00272_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12676_ net254 net2079 net432 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ net1220 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
X_11627_ _05880_ net660 vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15395_ clknet_leaf_27_wb_clk_i _01535_ _00203_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10034__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14346_ net1176 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XANTENNA__09975__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ net999 _07048_ net947 vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap316 _03596_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
Xhold608 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10509_ _06018_ _06019_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or3_1
XANTENNA__09196__Y _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold619 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ net1172 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
X_11489_ net655 _06356_ _06981_ _06982_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__o31a_1
XFILLER_0_12_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09188__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16016_ clknet_leaf_30_wb_clk_i _02156_ _00824_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13228_ net620 net936 net1021 net1451 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09727__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13159_ net232 _06991_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13287__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _03431_ _03436_ _03440_ _03441_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__a211o_1
XANTENNA__12495__A0 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _03336_ _03341_ _03361_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__and3_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ net2519 net1065 net35 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a21o_1
X_09321_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\] net711 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ _04837_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08716__B _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10273__A2 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] net898 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11470__B2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ _03917_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09183_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] net775 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09387__X _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ _03780_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09966__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08065_ _03782_ _03786_ _03755_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout1134_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09179__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_A _07192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16436__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] net743 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_A _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13278__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _03627_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nor2_1
X_08898_ net28 net1029 net986 net2352 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__o22a_1
XANTENNA__09351__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07849_ _03546_ net329 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10996__X _06508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10860_ _06373_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ net970 net631 net543 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _05314_ net386 vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12530_ net326 net2504 net447 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12461_ net312 net2622 net450 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14200_ net1184 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XANTENNA__10016__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _06205_ _06909_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__xnor2_1
X_15180_ net1140 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XANTENNA__09957__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net310 net2008 net459 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14131_ net1081 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11343_ _05294_ _05934_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14062_ net1075 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XANTENNA__09709__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ _05167_ net660 net657 _05168_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__a22o_1
X_13013_ _07452_ _07532_ _07453_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__o21a_1
X_10225_ team_02_WB.instance_to_wrap.top.a1.instruction\[24\] net791 net650 _05741_
+ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a22o_2
XANTENNA__15803__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\] net920 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a221o_1
XANTENNA__13269__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\] vssd1 vssd1 vccd1 vccd1
+ net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12103__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _05579_ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__nand2_1
X_14964_ net1238 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XANTENNA__09342__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16703_ net1345 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
X_13915_ net1261 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XANTENNA__11227__B _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14895_ net1221 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload3_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16634_ clknet_leaf_95_wb_clk_i _02753_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13426__C1 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13846_ net1147 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13777_ net2404 _03269_ net960 vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_187_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16565_ clknet_leaf_88_wb_clk_i _02689_ _01372_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13218__A1_N net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _04783_ _06028_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__xor2_1
XFILLER_0_186_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15516_ clknet_leaf_20_wb_clk_i _01656_ _00324_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10255__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12728_ _06841_ _06893_ _07251_ _06867_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__nor4b_1
XANTENNA__16309__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ clknet_leaf_127_wb_clk_i _02630_ _01303_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15447_ clknet_leaf_120_wb_clk_i _01587_ _00255_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12659_ net315 net1845 net435 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10007__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15378_ clknet_leaf_83_wb_clk_i _01518_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14329_ net1091 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
Xhold405 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] net757 net838 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a22o_1
Xfanout907 _04524_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_2
Xfanout918 _04515_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_55_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 _04511_ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09581__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ net2070 net1038 net990 team_02_WB.instance_to_wrap.ramaddr\[10\] vssd1 vssd1
+ vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
Xhold1105 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 team_02_WB.instance_to_wrap.top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1 net2478
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net847 _04360_ _04368_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__and3_1
Xhold1127 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12013__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09333__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07703_ _03392_ _03421_ _03390_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_178_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08683_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__or4_1
XANTENNA__11852__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07634_ team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] _03353_ team_02_WB.instance_to_wrap.top.a1.dataIn\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07631__A team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07565_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _03305_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_193_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout342_A _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13432__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _04814_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_192_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10246__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09235_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\] net673 _04748_ _04751_
+ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211o_1
XANTENNA__12683__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout607_A _06281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\] net815 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\]
+ _04674_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08117_ _03793_ _03830_ _03831_ _03790_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09097_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\] net753 net725 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08048_ _03765_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold950 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 team_02_WB.instance_to_wrap.top.a1.row1\[108\] vssd1 vssd1 vccd1 vccd1 net2323
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout976_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13808__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold983 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] net759 _05525_ _05526_
+ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__a211o_1
X_09999_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] net768 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ net312 net2459 net585 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_X clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11762__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _05956_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__or2_1
X_13700_ net1582 _03221_ net1066 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_103_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11682__A1 _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14680_ net1196 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
XANTENNA__07886__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net307 net2236 net488 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
XANTENNA__08637__A team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13631_ team_02_WB.instance_to_wrap.top.a1.row1\[101\] _03162_ vssd1 vssd1 vccd1
+ vccd1 _03181_ sky130_fd_sc_hd__and2_1
X_10843_ net414 net400 net545 vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11434__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13562_ net1050 _03113_ _03115_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__and4b_4
X_16350_ clknet_leaf_1_wb_clk_i _02490_ _01158_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07638__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10774_ net501 net385 vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_181_Right_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15301_ clknet_leaf_66_wb_clk_i _01445_ _00114_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12513_ net259 net2156 net446 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__mux2_1
X_16281_ clknet_leaf_123_wb_clk_i _02421_ _01089_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ _03061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.button_i
+ sky130_fd_sc_hd__inv_2
XANTENNA__12593__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ net236 net1937 net450 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__mux2_1
X_15232_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[23\]
+ _00045_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ net1157 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12375_ net641 _07195_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__nand2_4
XFILLER_0_62_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14114_ net1130 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
X_11326_ net421 _06037_ _06070_ _06104_ _06823_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__a32oi_2
X_15094_ net1078 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11937__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ net1203 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11257_ team_02_WB.instance_to_wrap.top.pc\[18\] _06263_ vssd1 vssd1 vccd1 vccd1
+ _06761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09563__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] net755 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a22o_1
X_11188_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__inv_2
XANTENNA__10173__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\] net730 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a22o_1
XANTENNA__13647__C1 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15996_ clknet_leaf_21_wb_clk_i _02136_ _00804_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09315__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14947_ net1137 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14878_ net1127 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12870__B1 _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16617_ clknet_leaf_90_wb_clk_i _02736_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13829_ net1155 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10228__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__B2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16548_ clknet_leaf_89_wb_clk_i _02672_ _01355_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16479_ clknet_leaf_83_wb_clk_i net1554 _01287_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08841__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09020_ net944 _04507_ _04509_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__and3_4
XFILLER_0_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11701__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15849__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold202 net186 vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold213 _02595_ vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_02_WB.instance_to_wrap.top.a1.hexop\[4\] vssd1 vssd1 vccd1 vccd1 net1586
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 team_02_WB.instance_to_wrap.top.a1.row2\[8\] vssd1 vssd1 vccd1 vccd1 net1597
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 _02606_ vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 team_02_WB.instance_to_wrap.ramstore\[10\] vssd1 vssd1 vccd1 vccd1 net1619
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11847__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold268 team_02_WB.instance_to_wrap.ramload\[27\] vssd1 vssd1 vccd1 vccd1 net1630
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\] vssd1
+ vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net781 _05434_ _05435_
+ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_1_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout704 _04389_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_4
XFILLER_0_111_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout715 _04385_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_8
Xfanout726 _04382_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
Xfanout737 _04379_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07626__A team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09853_ _05363_ _05365_ _05367_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4_1
Xfanout748 _04377_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_A _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net125 net1045 net992 net1472 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
X_09784_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\] net747 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a221o_1
XANTENNA__13638__C1 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08735_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\] net932 team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__and3b_2
XANTENNA__12678__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_1_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07617_ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1 vccd1 _03340_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08597_ _04254_ _04255_ _04256_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout724_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11416__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1
+ _03289_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08744__X _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09218_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10490_ _05559_ _06006_ net510 _05556_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_20_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__A1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] net751 _04664_ _04665_
+ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14922__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12160_ net302 net2619 net465 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
XANTENNA__09793__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11757__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _06230_ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__xnor2_1
X_12091_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] net292 net581 vssd1
+ vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
Xhold780 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net667 _06541_ _06548_ net656 vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__o22a_1
XANTENNA__08899__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ clknet_leaf_32_wb_clk_i _01990_ _00658_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16154__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14801_ net1231 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15781_ clknet_leaf_26_wb_clk_i _01921_ _00589_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12993_ _07475_ _07512_ _07473_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14732_ net1215 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11944_ net236 net2373 net584 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11875_ net244 net2360 net487 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15261__Q team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14663_ net1181 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16402_ clknet_leaf_100_wb_clk_i _02537_ _01210_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_10826_ _06335_ _06341_ net394 vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__mux2_1
X_13614_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] _03108_ vssd1 vssd1 vccd1
+ vccd1 _03166_ sky130_fd_sc_hd__nor2_1
XANTENNA__11407__B2 _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09076__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14594_ net1130 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16333_ clknet_leaf_51_wb_clk_i _02473_ _01141_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13545_ _03080_ _03101_ _03102_ net1068 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__o211a_1
X_10757_ net999 _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nor2_1
XANTENNA__08823__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13476_ team_02_WB.START_ADDR_VAL_REG\[16\] net1071 net1005 vssd1 vssd1 vccd1 vccd1
+ net199 sky130_fd_sc_hd__a21o_1
X_16264_ clknet_leaf_24_wb_clk_i _02404_ _01072_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ net789 _04419_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__o21a_2
X_12427_ net304 net2376 net457 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
X_15215_ clknet_leaf_98_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[6\]
+ _00028_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12907__B2 _05017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16195_ clknet_leaf_9_wb_clk_i _02335_ _01003_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09784__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ net300 net2148 net562 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
X_15146_ net1144 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11309_ _06262_ _06810_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__or2_1
XANTENNA_max_cap522_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15077_ net1246 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
X_12289_ net272 net2226 net570 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
X_14028_ net1215 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_0__f_wb_clk_i_X clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire525_A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15979_ clknet_leaf_15_wb_clk_i _02119_ _00787_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11255__X _06759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\] net979 vssd1 vssd1 vccd1
+ vccd1 _04209_ sky130_fd_sc_hd__or2_1
XANTENNA__10600__A _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08451_ _04145_ _04153_ _04148_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__or3b_1
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08382_ _04059_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09067__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15671__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08814__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10082__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09003_ _04510_ _04519_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__nor2_4
XFILLER_0_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout305_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13358__A net2158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1214_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13049__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\] net725 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\]
+ _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 _07223_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_8
Xfanout567 _07218_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_4
X_09836_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\] net766 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__a22o_1
Xfanout578 _07214_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_6
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_198_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout841_A _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _05277_ _05279_ _05281_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or4_1
XANTENNA__14189__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12201__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ _04268_ _04346_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__nor2_4
X_09698_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\] net726 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_202_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08649_ net1061 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11660_ _05738_ _05916_ _07141_ _07145_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__or4b_1
XFILLER_0_138_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09058__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10611_ _04283_ _04493_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__nand2_8
XFILLER_0_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ net670 _07075_ _07079_ net836 vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10073__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ team_02_WB.instance_to_wrap.top.a1.hexop\[1\] team_02_WB.instance_to_wrap.top.a1.hexop\[2\]
+ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__or3_1
X_10542_ net389 _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13261_ net1462 net983 net965 _02978_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ net519 _05333_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__nand2_1
X_12212_ net2136 net245 net615 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__mux2_1
X_15000_ net1133 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
XANTENNA__09766__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13192_ _07390_ _07392_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09230__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08650__A team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12143_ _06278_ _07190_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__nor2_2
XANTENNA__13268__A _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13314__B2 _03006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ net350 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] net470 vssd1
+ vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
XANTENNA__11325__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _06534_ _06535_ net412 vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__mux2_1
X_15902_ clknet_leaf_5_wb_clk_i _02042_ _00710_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15833_ clknet_leaf_124_wb_clk_i _01973_ _00641_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15764_ clknet_leaf_114_wb_clk_i _01904_ _00572_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12111__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ team_02_WB.instance_to_wrap.top.pc\[2\] _05835_ vssd1 vssd1 vccd1 vccd1 _07496_
+ sky130_fd_sc_hd__xnor2_1
X_14715_ net1077 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
X_11927_ net314 net2022 net484 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
X_15695_ clknet_leaf_48_wb_clk_i _01835_ _00503_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11950__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14827__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14646_ net1120 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
X_11858_ net307 net2367 net493 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ _04755_ net405 vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_171_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14577_ net1229 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11789_ net297 net1892 net594 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ clknet_leaf_20_wb_clk_i _02456_ _01124_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10603__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _03084_ _03085_ _03087_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__or4_1
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16247_ clknet_leaf_122_wb_clk_i _02387_ _01055_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09927__Y _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ team_02_WB.START_ADDR_VAL_REG\[0\] _03309_ net1003 vssd1 vssd1 vccd1 vccd1
+ _03060_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09757__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
X_16178_ clknet_leaf_76_wb_clk_i _02318_ _00986_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09221__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__13178__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15129_ net1158 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09509__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _03670_ _03672_ _03660_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13305__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13906__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _03585_ _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_182_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09391__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] net750 net714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a22o_1
X_09552_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\] net909 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a22o_1
XANTENNA__11619__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12816__B1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ team_02_WB.instance_to_wrap.top.a1.data\[8\] net958 _04196_ vssd1 vssd1 vccd1
+ vccd1 _04197_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09483_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\] net682 _04998_ _04999_
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout255_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ _04127_ _04133_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08365_ _04041_ _04054_ _04074_ _04053_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout422_A _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08296_ _03962_ _03988_ _03985_ _03980_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__a211o_1
XANTENNA__09460__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12691__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09748__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1158_X net2520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_86_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout320 _06936_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_167_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout331 _07013_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_1
Xfanout342 _07051_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
Xfanout353 _07126_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_204_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout364 _07107_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_2
Xfanout375 _06088_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_2
Xfanout386 _05901_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_2
XANTENNA__09920__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout397 net400 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_4
X_09819_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _04588_ _06130_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__nor2_1
XANTENNA__09279__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12761_ _04823_ _04909_ _05083_ _05168_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__or4_1
XANTENNA__11770__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10294__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14500_ net1100 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ net262 net1796 net603 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15480_ clknet_leaf_123_wb_clk_i _01620_ _00288_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12692_ net314 net1849 net432 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11643_ _05995_ _06287_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14431_ net1115 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
XANTENNA__13232__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09987__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11574_ _06583_ _07059_ _07060_ _07063_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__o211ai_2
X_14362_ net1096 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11794__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16101_ clknet_leaf_29_wb_clk_i _02241_ _00909_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10525_ _05877_ net402 vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__nor2_1
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13313_ team_02_WB.instance_to_wrap.top.pc\[3\] net1056 _07083_ net934 vssd1 vssd1
+ vccd1 vccd1 _03006_ sky130_fd_sc_hd__a22o_1
X_14293_ net1257 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XANTENNA__08651__Y _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09476__A _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16032_ clknet_leaf_17_wb_clk_i _02172_ _00840_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09739__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ _06415_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_1
X_10456_ _05080_ _05061_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09203__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13175_ net1026 _02936_ net1023 team_02_WB.instance_to_wrap.top.pc\[6\] vssd1 vssd1
+ vccd1 vccd1 _01487_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10415__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__inv_2
XANTENNA__12106__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ net300 net2388 net467 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XANTENNA__11945__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ net284 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\] net470 vssd1
+ vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
X_11008_ _04777_ net661 net659 _04782_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09911__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15816_ clknet_leaf_25_wb_clk_i _01956_ _00624_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_16796_ net1340 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15747_ clknet_leaf_8_wb_clk_i _01887_ _00555_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12959_ team_02_WB.instance_to_wrap.top.pc\[11\] _05444_ vssd1 vssd1 vccd1 vccd1
+ _07479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10285__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ clknet_leaf_5_wb_clk_i _01818_ _00486_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14629_ net1114 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13223__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ _03796_ _03824_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09978__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09442__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__A0 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08081_ _03774_ net228 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__xor2_2
XFILLER_0_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14292__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11537__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12016__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ net1058 net952 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and2_1
XANTENNA__11855__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13636__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07934_ _03608_ _03653_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_149_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09902__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ _03556_ _03586_ _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout372_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _05107_ _05115_ _05118_ _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__nor4_1
XFILLER_0_97_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ _03490_ _03497_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__o21a_1
XFILLER_0_211_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\] net759 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12686__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout637_A _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10276__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13371__A net2397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09466_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\] net828 net866 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_195_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08465__A team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08417_ _04113_ _04122_ _04124_ _04109_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o2bb2a_2
X_09397_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] net754 net711 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\]
+ _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a221o_1
XANTENNA__13214__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_A _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10028__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04059_ vssd1 vssd1 vccd1
+ vccd1 _04060_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10579__A1 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08752__X _04381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08279_ _03962_ _03988_ _03976_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1
+ vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10310_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\] net781 _05818_ _05819_
+ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11290_ _05212_ _06016_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_91_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10241_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] net822 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\]
+ _05744_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10200__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _05673_ _05684_ _05686_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__nor4_1
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__buf_4
Xfanout1115 net1118 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_4
XANTENNA__11765__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1128 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_4
Xfanout1137 net1138 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__buf_4
X_14980_ net1156 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1148 net1149 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_2
Xfanout1159 net1161 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_2
X_13931_ net1259 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11700__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16650_ clknet_leaf_94_wb_clk_i _02769_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13862_ net1149 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15601_ clknet_leaf_0_wb_clk_i _01741_ _00409_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12813_ team_02_WB.instance_to_wrap.top.testpc.en_latched team_02_WB.instance_to_wrap.top.i_ready
+ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__and2_2
X_16581_ clknet_leaf_92_wb_clk_i _02700_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12596__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13793_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ _03278_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15532_ clknet_leaf_2_wb_clk_i _01672_ _00340_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12744_ _06667_ _06700_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_177_Left_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09672__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ clknet_leaf_42_wb_clk_i _01603_ _00271_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13205__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12675_ net237 net1909 net430 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14414_ net1076 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _05902_ _05996_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15394_ clknet_leaf_116_wb_clk_i _01534_ _00202_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14345_ net1221 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
Xwire540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11557_ _06255_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10508_ _06022_ _06024_ _05984_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
X_11488_ _06977_ _06981_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__or2_1
X_14276_ net1099 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16015_ clknet_leaf_43_wb_clk_i _02155_ _00823_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10439_ _04695_ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__nor2_1
X_13227_ net621 net937 net1022 net1394 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_186_Left_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ net1026 _02922_ net1023 team_02_WB.instance_to_wrap.top.pc\[9\] vssd1 vssd1
+ vccd1 vccd1 _01490_ sky130_fd_sc_hd__a2bb2o_1
X_12109_ _06278_ _07188_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nor2_1
X_13089_ _06707_ net234 net231 _02863_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11298__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13692__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07650_ _03336_ _03361_ _03341_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_195_Right_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07581_ net2407 net1065 net36 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a21o_1
X_16779_ net1323 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
X_09320_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] net768 net744 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a22o_1
XANTENNA__10258__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\] net816 net804 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\]
+ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08871__B1 _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08202_ _03884_ _03918_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] net754 net706 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\]
+ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09415__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ _03842_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_190_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10607__X _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _03706_ _03784_ _03785_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__nor3_2
XFILLER_0_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1127_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11930__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13366__A team_02_WB.instance_to_wrap.ramload\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08966_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\] net695 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a22o_1
XANTENNA__15605__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ _03571_ _03600_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and2_1
XANTENNA__10061__Y _05578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13683__B1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net29 net1032 net988 net2568 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout754_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ _03537_ _03569_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__xor2_2
XANTENNA__08747__X _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15755__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14197__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10249__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ _05020_ _05021_ _05030_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__nor4_2
XFILLER_0_94_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10790_ _06304_ _06305_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__or2_1
XANTENNA__11997__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09449_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\] net757 _04964_ _04965_
+ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08862__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13232__A2_N net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ net305 net2118 net452 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09406__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__A team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08614__A0 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11411_ _03294_ net848 vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__or2_1
X_12391_ net303 net2383 net460 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ net670 _06841_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__nand2_1
X_14130_ net1183 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_115_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11273_ _06546_ _06773_ net413 vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__mux2_1
X_14061_ net1121 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input50_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _05693_ _05740_ net550 vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__mux2_1
X_13012_ team_02_WB.instance_to_wrap.top.pc\[25\] _06172_ _07531_ vssd1 vssd1 vccd1
+ vccd1 _07532_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09754__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] net822 net908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15285__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14963_ net1079 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
Xhold6 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\] vssd1 vssd1 vccd1 vccd1
+ net1368 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _05583_ _05602_ net968 vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__mux2_1
XANTENNA__15264__Q team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16702_ net1344 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_13914_ net1229 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14894_ net1076 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XANTENNA__09893__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16633_ clknet_leaf_95_wb_clk_i _02752_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13845_ net1151 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11437__C1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16564_ clknet_leaf_88_wb_clk_i _02688_ _01371_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13776_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] _03269_
+ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__and2_1
X_10988_ _05954_ _06499_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09645__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15515_ clknet_leaf_34_wb_clk_i _01655_ _00323_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12727_ _06957_ _07250_ _06915_ _06937_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16495_ clknet_leaf_0_wb_clk_i _02629_ _01302_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08853__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15446_ clknet_leaf_50_wb_clk_i _01586_ _00254_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12658_ net306 net2553 net437 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08605__A0 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ _05833_ _05998_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15377_ clknet_leaf_83_wb_clk_i _01517_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12589_ net302 net2585 net441 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14328_ net1195 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_194_Left_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold406 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold417 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14259_ net1072 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08908__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08908__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09030__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 _04524_ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 _04515_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_55_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ net1587 net1038 net990 team_02_WB.instance_to_wrap.ramaddr\[11\] vssd1 vssd1
+ vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XANTENNA__10191__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ net846 _04368_ _04370_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__and3_4
Xhold1128 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1139 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
X_07702_ _03422_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__nor2_1
XANTENNA__09670__Y _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08682_ net1062 _04308_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand2_1
XANTENNA__11140__A1 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09884__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07633_ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] _03339_ _03342_ _03344_ _03355_
+ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__o41a_2
X_07564_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 _03304_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09097__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09636__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09303_ _04816_ _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__or3_1
XANTENNA__08844__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout335_A _06994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1077_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13028__B1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\] net741 _04749_ _04750_
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09839__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\] net830 net925 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\]
+ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1244_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ _03832_ _03834_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\] net733 net705 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08047_ _03725_ _03752_ _03767_ _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold940 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold951 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_A _04496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12204__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] net752 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a22o_1
XANTENNA__10182__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ _04270_ _04273_ _04457_ _04465_ _04309_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13120__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ net304 net2368 net587 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_1
XANTENNA__09875__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _04695_ _05955_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__and2_1
X_11891_ net299 net1530 net487 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13630_ net1411 net962 _03180_ net1067 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__o211a_1
X_10842_ net545 net419 vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__and2_1
XANTENNA__09088__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ _03289_ net1049 _03113_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__and4_1
XANTENNA__08835__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ net608 net402 vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15300_ clknet_leaf_70_wb_clk_i _01444_ _00113_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12512_ net250 net2113 net448 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16280_ clknet_leaf_123_wb_clk_i _02420_ _01088_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce_dly team_02_WB.instance_to_wrap.top.pad.button_control.debounce
+ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and2b_4
XANTENNA_input98_A wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[22\]
+ _00044_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\]
+ sky130_fd_sc_hd__dfrtp_2
X_12443_ net244 net2128 net452 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ net1157 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
X_12374_ net347 net2084 net560 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14113_ net1261 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
X_11325_ _05988_ net664 net656 _06825_ _06824_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_97_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15093_ net1080 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
X_11256_ _06218_ _06219_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__xnor2_1
X_14044_ net1192 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09563__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\] net744 net716 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a22o_1
XANTENNA__11519__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ net410 _06449_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12114__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10138_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] net782 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\]
+ _05654_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15995_ clknet_leaf_32_wb_clk_i _02135_ _00803_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11953__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13293__X _02996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\] net917 net873 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a22o_1
X_14946_ net1129 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
XANTENNA__09866__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14877_ net1203 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16616_ clknet_leaf_90_wb_clk_i _02735_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09079__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ net1149 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09618__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16547_ clknet_leaf_89_wb_clk_i _02671_ _01354_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_13759_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or2_1
XANTENNA__15300__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16478_ clknet_leaf_83_wb_clk_i net1559 _01286_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15429_ clknet_leaf_29_wb_clk_i _01569_ _00237_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09251__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 team_02_WB.instance_to_wrap.ramstore\[3\] vssd1 vssd1 vccd1 vccd1 net1576
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13909__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold225 net108 vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 team_02_WB.instance_to_wrap.top.a1.row1\[3\] vssd1 vssd1 vccd1 vccd1 net1609
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_02_WB.instance_to_wrap.top.a1.hexop\[2\] vssd1 vssd1 vccd1 vccd1 net1620
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\] net773 _05436_ _05437_
+ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__a211o_1
Xhold269 team_02_WB.instance_to_wrap.ramaddr\[13\] vssd1 vssd1 vccd1 vccd1 net1631
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 net708 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_8
Xfanout716 _04385_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_4
X_09852_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\] net828 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a221o_1
Xfanout727 _04382_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12024__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout738 _04379_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
Xfanout749 net750 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10164__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ net126 net1045 net992 net1462 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
X_09783_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] net776 net704 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11863__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A _06766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__and3b_2
XANTENNA__08738__A team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13363__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _03298_ _04278_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1194_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07616_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03338_ vssd1 vssd1 vccd1
+ vccd1 _03339_ sky130_fd_sc_hd__xnor2_1
X_08596_ net56 net55 net58 net57 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__or4_4
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12694__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11416__A2 _06908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08817__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout717_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09490__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _04714_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12916__A2 _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__A1_N net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\] net775 net767 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a22o_1
XANTENNA__09242__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__X _04389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] net887 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13819__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12129__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15943__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11110_ _06174_ _06175_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net1651 net284 net580 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
Xhold770 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold781 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13217__A1_N _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ net382 _06104_ _06549_ _06531_ _06110_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a32o_1
Xhold792 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10155__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ net1260 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15780_ clknet_leaf_34_wb_clk_i _01920_ _00588_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12992_ _07476_ _07511_ _07477_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09848__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14731_ net1152 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ net247 net2211 net586 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ net1205 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ net241 net1563 net487 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
X_16401_ clknet_leaf_88_wb_clk_i _02536_ _01209_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13613_ net1049 _03114_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11407__A2 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ _06337_ _06340_ net369 vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08808__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14593_ net1259 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16332_ clknet_leaf_2_wb_clk_i _02472_ _01140_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13544_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] _03061_ vssd1 vssd1 vccd1
+ vccd1 _03102_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09481__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10756_ team_02_WB.instance_to_wrap.top.pc\[31\] _06272_ vssd1 vssd1 vccd1 vccd1
+ _06273_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16263_ clknet_leaf_39_wb_clk_i _02403_ _01071_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ team_02_WB.START_ADDR_VAL_REG\[15\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net198 sky130_fd_sc_hd__a21o_1
X_10687_ net994 net550 _04417_ _06127_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a31o_1
XFILLER_0_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15214_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[5\]
+ _00027_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ net297 net1936 net456 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__mux2_1
X_16194_ clknet_leaf_102_wb_clk_i _02334_ _01002_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11948__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ net1158 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12357_ net294 net1758 net561 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11591__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11308_ team_02_WB.instance_to_wrap.top.pc\[15\] _06261_ team_02_WB.instance_to_wrap.top.pc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__a21oi_1
X_15076_ net1245 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
X_12288_ net289 net1965 net569 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
X_14027_ net1124 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
X_11239_ net668 _06742_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10146__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13464__A team_02_WB.START_ADDR_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15978_ clknet_leaf_38_wb_clk_i _02118_ _00786_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13096__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__X _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14929_ net1231 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XFILLER_0_210_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08450_ _04145_ _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04070_ vssd1 vssd1 vccd1
+ vccd1 _04091_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_175_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09389__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12019__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09002_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ net1058 net952 vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o31a_2
XANTENNA__09224__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11858__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09904_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] net741 net685 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1148_A team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10137__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1207_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 _04489_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout557 _07223_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
X_09835_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] net778 net698 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\]
+ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a221o_1
Xfanout568 _07217_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12689__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 _07214_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_4
XANTENNA__11446__X _06942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] net928 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a221o_1
X_08717_ _04288_ _04320_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nand2_2
XANTENNA__11606__B _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\] net745 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout834_A _04506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10845__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08648_ _03298_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04277_ sky130_fd_sc_hd__or2_2
XFILLER_0_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ net1724 _04241_ _04225_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10610_ _04283_ _04493_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__and2_2
XFILLER_0_181_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11590_ _05906_ _05910_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08634__C team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net517 net386 _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_134_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ team_02_WB.instance_to_wrap.top.pc\[28\] net1055 net934 _02977_ vssd1 vssd1
+ vccd1 vccd1 _02978_ sky130_fd_sc_hd__a22o_1
X_10472_ _05295_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11768__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ net2009 net241 net614 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ _07334_ _07496_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11573__A1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11573__B2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ net346 net2214 net466 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
XANTENNA__13268__B _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12073_ net362 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\] net470 vssd1
+ vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
X_11024_ _06381_ _06384_ net395 vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__mux2_1
X_15901_ clknet_leaf_10_wb_clk_i _02041_ _00709_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12599__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ clknet_leaf_114_wb_clk_i _01972_ _00640_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13078__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ clknet_leaf_47_wb_clk_i _01903_ _00571_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11628__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15272__Q team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ _07493_ _07494_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14714_ net1087 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
X_11926_ net306 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\] net485 vssd1
+ vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15694_ clknet_leaf_45_wb_clk_i _01834_ _00502_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10300__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14645_ net1242 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
X_11857_ net296 net2481 net492 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15989__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10808_ _04802_ net387 vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nor2_1
X_14576_ net1234 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ net311 net2475 net593 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16315_ clknet_leaf_34_wb_clk_i _02455_ _01123_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13527_ _03081_ _03082_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__nor2_1
X_10739_ team_02_WB.instance_to_wrap.top.pc\[7\] team_02_WB.instance_to_wrap.top.pc\[6\]
+ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16246_ clknet_leaf_50_wb_clk_i _02386_ _01054_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13458_ _02768_ _03047_ _03059_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09206__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12409_ net242 net1766 net456 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
X_16177_ clknet_leaf_1_wb_clk_i _02317_ _00985_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13389_ team_02_WB.instance_to_wrap.ramload\[18\] net1011 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[18\] sky130_fd_sc_hd__and2_1
XFILLER_0_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10367__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
X_15128_ net1158 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10154__Y _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15369__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13305__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _03670_ _03672_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__and2_1
X_15059_ net1251 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XANTENNA__10119__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ net316 _03597_ _03581_ _03584_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a211o_1
XFILLER_0_207_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09620_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] net730 _05134_ _05136_
+ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a211o_1
XANTENNA__12302__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\] net826 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ _05067_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a221o_1
XANTENNA__11619__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08502_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\] net979 vssd1 vssd1 vccd1
+ vccd1 _04196_ sky130_fd_sc_hd__or2_1
XFILLER_0_195_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09482_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] net709 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08433_ _04128_ _04130_ _04133_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout248_A _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08364_ _04030_ _04053_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nand3_1
XFILLER_0_160_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14753__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ _03962_ _03988_ _03980_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13529__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16144__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1265_A team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11555__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__B team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08971__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout310 _06840_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout321 _06955_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_2
Xfanout332 _07013_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_2
Xfanout343 _07051_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_1
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 net357 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_204_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout365 _07107_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_1
Xfanout376 net377 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_2
X_09818_ _05314_ _05333_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or2_1
Xfanout398 net399 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12212__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09749_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] net771 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ _04694_ _05252_ _05335_ _05420_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11711_ net268 net1525 net602 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XANTENNA__11491__B1 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ net305 net2234 net433 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11352__A _06104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14430_ net1128 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
X_11642_ net547 net385 vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09436__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14361_ net1097 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11573_ net836 _07057_ _07058_ net668 _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16100_ clknet_leaf_34_wb_clk_i _02240_ _00908_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_13312_ net1584 net984 net967 _03005_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input80_A wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10524_ _06039_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or2_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_1
X_14292_ net1153 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
X_16031_ clknet_leaf_61_wb_clk_i _02171_ _00839_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13243_ _06458_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__nor2_1
X_10455_ _05061_ _05080_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__and2b_1
XANTENNA__10349__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13174_ _07027_ net232 _02933_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__o211a_1
X_10386_ _05880_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15267__Q team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ net294 net1725 net468 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
XANTENNA__08962__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_176_Right_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13299__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ net273 net2607 net472 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _04783_ net664 _06410_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12122__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15815_ clknet_leaf_41_wb_clk_i _01955_ _00623_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_16795_ net1339 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__11961__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15746_ clknet_leaf_119_wb_clk_i _01886_ _00554_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12958_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__inv_2
XANTENNA__09675__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ net244 net2188 net484 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15677_ clknet_leaf_4_wb_clk_i _01817_ _00485_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12889_ _07407_ _07408_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16167__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14628_ net1099 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XANTENNA__09003__Y _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13223__B2 _05510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14559_ net1116 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XANTENNA__14573__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08080_ _03795_ _03800_ _03790_ _03792_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16229_ clknet_leaf_28_wb_clk_i _02369_ _01037_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__C1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08982_ net997 _04310_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__or2_1
XANTENNA_wire540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__inv_2
XANTENNA__08510__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09902__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _03571_ _03574_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__nand2b_2
XANTENNA__12032__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09603_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\] net809 net869 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\]
+ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ _03465_ _03474_ net366 _03488_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout365_A _07107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14748__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09534_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] net779 net735 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09666__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13371__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09130__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\] _04981_ vssd1 vssd1 vccd1
+ vccd1 _04982_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08416_ _04104_ _04115_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09396_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] net771 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__a22o_1
XANTENNA__09418__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08347_ _04047_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_102_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08278_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] _03989_ vssd1 vssd1 vccd1
+ vccd1 _03993_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_78_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout999_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12207__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10240_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\] net908 _05743_ _05756_
+ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_91_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10171_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] net834 net915 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\]
+ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a221o_1
Xfanout1105 net1110 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1116 net1118 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_2
Xfanout1127 net1128 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_4
XFILLER_0_206_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1138 net1171 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_4
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1151 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_4
X_13930_ net1259 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_98_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11700__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13861_ net1151 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11781__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15600_ clknet_leaf_30_wb_clk_i _01740_ _00408_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12812_ net231 _07334_ _07335_ _07329_ _04280_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a32o_1
X_16580_ clknet_leaf_91_wb_clk_i _02699_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dfxtp_1
X_13792_ _03280_ _03281_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09657__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09121__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15531_ clknet_leaf_15_wb_clk_i _01671_ _00339_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12743_ _06728_ _06754_ _07266_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__nand3_1
XFILLER_0_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10267__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ clknet_leaf_7_wb_clk_i _01602_ _00270_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12674_ net245 net1976 net432 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08880__B2 net2520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10019__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14413_ net1126 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
X_11625_ net421 _06776_ _07111_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__o21a_1
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ clknet_leaf_103_wb_clk_i _01533_ _00201_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_X clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ net1113 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire541 _04754_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11556_ team_02_WB.instance_to_wrap.top.pc\[5\] _06254_ vssd1 vssd1 vccd1 vccd1 _07047_
+ sky130_fd_sc_hd__nor2_1
X_10507_ _05972_ _05976_ _06023_ _06020_ _05977_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o32a_1
XFILLER_0_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14275_ net1137 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XANTENNA__12117__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11487_ net376 _06796_ _06980_ net383 vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__a22o_1
X_16014_ clknet_leaf_46_wb_clk_i _02154_ _00822_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13226_ net646 net936 net1021 net1383 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09188__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10438_ _04779_ _05954_ _04734_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11956__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ _06972_ net232 _02921_ net976 _02919_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__o221a_1
X_10369_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\] net874 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12108_ net1962 net347 net580 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
X_13088_ _07365_ _07426_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__xnor2_1
X_12039_ net363 net2215 net474 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09896__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ net2111 net1065 net37 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a21o_1
X_16778_ net1322 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XANTENNA__09648__B1 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09112__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09014__X _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15729_ clknet_leaf_126_wb_clk_i _01869_ _00537_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] net926 net910 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_177_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08871__A1 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ _03886_ _03898_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__xor2_2
X_09181_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\] net782 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08132_ _03850_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_190_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09820__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ _03711_ _03753_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12027__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09179__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11866__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1022_A _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__C1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13366__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\] net746 _04473_ _04475_
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a2111o_2
XANTENNA_fanout482_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _03605_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and2_1
XANTENNA__09887__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ net30 net1029 net986 net2249 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__o22a_1
XANTENNA__09351__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__A _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _03537_ _03551_ net329 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_197_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_X clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07778_ _03467_ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09103__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] net866 _05031_ _05033_
+ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a211o_1
X_16755__1299 vssd1 vssd1 vccd1 vccd1 _16755__1299/HI net1299 sky130_fd_sc_hd__conb_1
XFILLER_0_211_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout914_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09448_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\] net785 net753 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09379_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] net807 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\]
+ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11410_ net670 _06893_ _06907_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_136_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12390_ net294 net2107 net460 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11341_ _05294_ _06015_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14060_ net1215 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11272_ net417 _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__nor2_1
XANTENNA__11776__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _07530_ _07454_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__and2b_1
X_10223_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] net648 _05739_ vssd1
+ vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a21o_1
XANTENNA__10185__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] net791 _05670_ vssd1
+ vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a21oi_4
X_14962_ net1177 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
X_10085_ _05594_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__or2_4
Xhold7 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\] vssd1 vssd1 vccd1 vccd1
+ net1369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09878__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ net1343 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_13913_ net1233 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14893_ net1120 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XANTENNA__14388__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08657__Y _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16632_ clknet_leaf_95_wb_clk_i _02751_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13844_ net1147 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
XANTENNA__12400__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13775_ _03269_ _03270_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__nor2_1
X_16563_ clknet_leaf_88_wb_clk_i _02687_ _01370_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ _04783_ _05953_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _06976_ _07014_ _07249_ _06995_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__and4bb_1
X_15514_ clknet_leaf_52_wb_clk_i _01654_ _00322_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16494_ clknet_leaf_0_wb_clk_i _02628_ _01301_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15445_ clknet_leaf_32_wb_clk_i _01585_ _00253_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12657_ net298 net1938 net436 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ net794 _07094_ _06117_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__o21a_1
X_15376_ clknet_leaf_83_wb_clk_i _01516_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__09802__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ net293 net2212 net439 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__mux2_1
XANTENNA__10948__C1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14327_ net1208 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
X_11539_ net1692 net338 net637 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XANTENNA__14851__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold407 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold429 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ net1183 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
X_13209_ net1453 net1021 net939 _04904_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14189_ net1128 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout909 _04524_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09009__X _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1107 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ net846 _04360_ _04365_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_146_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1118 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1129 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ _03383_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__xor2_1
XANTENNA__09333__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08681_ net1063 net1062 _04266_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_179_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07632_ _03328_ _03346_ _03352_ team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] team_02_WB.instance_to_wrap.top.a1.dataIn\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_178_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12310__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07563_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_76_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\] net900 net797 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ _04808_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09233_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\] net781 net745 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] net908 net895 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08115_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_211_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09095_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\] net677 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10066__A _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1237_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _03744_ _03750_ _03766_ _03725_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_170_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold930 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold941 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold952 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13377__A net2411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09572__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _05489_ _05511_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _04310_ _04316_ _04317_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__nand3_1
X_08879_ net17 net1029 net986 net2514 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10910_ net2134 net239 net638 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XANTENNA__12220__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ net310 net2608 net489 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15872__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _06355_ _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nand2_2
XFILLER_0_168_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__nor2_2
X_10772_ _06286_ _06287_ net390 vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12511_ net253 net2356 net448 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__mux2_1
XANTENNA__10642__A1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ team_02_WB.START_ADDR_VAL_REG\[31\] net1071 net1004 vssd1 vssd1 vccd1 vccd1
+ net216 sky130_fd_sc_hd__a21o_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15230_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[21\]
+ _00043_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_117_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ net240 net2600 net453 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15161_ net1144 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
X_12373_ net350 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\] net560 vssd1
+ vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14112_ net1102 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
X_11324_ _06358_ _06821_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__or2_1
X_15092_ net1074 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
X_14043_ net1075 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
X_11255_ _06743_ _06756_ _06758_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__or3b_4
XPHY_EDGE_ROW_26_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10158__B1 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__Y _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] net783 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\]
+ _05722_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a221o_1
XANTENNA__09563__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ net409 _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\] net746 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15994_ clknet_leaf_19_wb_clk_i _02134_ _00802_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09315__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14945_ net1256 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\] net808 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15007__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10330__B1 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14876_ net1193 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16615_ clknet_leaf_90_wb_clk_i _02734_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13827_ net1149 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13758_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__nand2_1
X_16546_ clknet_leaf_88_wb_clk_i _02670_ _01353_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_190_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12709_ net848 _04355_ _06162_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13689_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\]
+ _03200_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16477_ clknet_leaf_83_wb_clk_i net1507 _01285_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13293__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15428_ clknet_leaf_36_wb_clk_i _01568_ _00236_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16721__1353 vssd1 vssd1 vccd1 vccd1 net1353 _16721__1353/LO sky130_fd_sc_hd__conb_1
XANTENNA_wire498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09946__Y _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15359_ clknet_leaf_73_wb_clk_i _01499_ _00172_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_170_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14581__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold204 team_02_WB.START_ADDR_VAL_REG\[23\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold215 team_02_WB.instance_to_wrap.top.a1.row1\[109\] vssd1 vssd1 vccd1 vccd1 net1577
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold226 _02605_ vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_02_WB.instance_to_wrap.top.a1.row1\[122\] vssd1 vssd1 vccd1 vccd1 net1599
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\] net701 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a22o_1
Xhold248 team_02_WB.instance_to_wrap.ramaddr\[22\] vssd1 vssd1 vccd1 vccd1 net1610
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 team_02_WB.instance_to_wrap.top.a1.row1\[10\] vssd1 vssd1 vccd1 vccd1 net1621
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10149__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12305__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16754__1298 vssd1 vssd1 vccd1 vccd1 _16754__1298/HI net1298 sky130_fd_sc_hd__conb_1
XANTENNA__10614__A _06130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net708 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout717 net720 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_8
X_09851_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\] net833 net821 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a22o_1
Xfanout728 _04382_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
Xfanout739 _04379_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_8
X_08802_ net127 net1045 net992 net1431 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
X_09782_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\] net759 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\]
+ _05296_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15895__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ net847 _04360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__and3_4
XFILLER_0_147_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12040__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _04291_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10321__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _03324_ _03328_ _03325_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__a21oi_1
X_08595_ net63 net62 net59 net60 vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__or4bb_4
XANTENNA_fanout445_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1187_A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ net971 net634 net544 vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09147_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] net783 net758 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14491__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_X net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09793__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\] net834 net928 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\]
+ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__X _06686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08029_ _03744_ _03750_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nand2_2
XANTENNA__12215__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold760 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\] vssd1
+ vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold782 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _05951_ net661 net658 _04823_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__a22o_1
XANTENNA__09545__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold793 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12991_ team_02_WB.instance_to_wrap.top.pc\[11\] _05445_ _07510_ vssd1 vssd1 vccd1
+ vccd1 _07511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_207_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14730_ net1117 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
X_11942_ net240 net2165 net586 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14661_ net1172 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ net643 _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12065__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16400_ clknet_leaf_100_wb_clk_i _02535_ _01208_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_13612_ _03160_ _03163_ _03108_ _03135_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _06338_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__or2_1
X_14592_ net1106 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16331_ clknet_leaf_16_wb_clk_i _02471_ _01139_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13543_ team_02_WB.instance_to_wrap.top.edg2.button_i _03090_ _03099_ _03100_ vssd1
+ vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__or4_1
XFILLER_0_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10755_ team_02_WB.instance_to_wrap.top.pc\[30\] _06271_ vssd1 vssd1 vccd1 vccd1
+ _06272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10091__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16262_ clknet_leaf_10_wb_clk_i _02402_ _01070_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13474_ team_02_WB.START_ADDR_VAL_REG\[14\] _04260_ vssd1 vssd1 vccd1 vccd1 net197
+ sky130_fd_sc_hd__and2_1
XFILLER_0_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_80_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10686_ _06201_ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15213_ clknet_leaf_97_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[4\]
+ _00026_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] sky130_fd_sc_hd__dfrtp_4
X_12425_ net308 net2115 net455 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
X_16193_ clknet_leaf_102_wb_clk_i _02333_ _01001_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10379__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144_ net1143 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XANTENNA__09784__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12356_ net284 net2509 net563 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__mux2_1
XANTENNA__08603__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13317__B1 _07122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _06214_ _06808_ net973 vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15075_ net1251 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XANTENNA__10434__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ net279 net2628 net568 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XANTENNA__12125__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ net1117 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XANTENNA__09536__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _05127_ _06597_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_52_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11964__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _06355_ _06674_ net656 vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__a21o_1
XANTENNA__07743__A team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13464__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15977_ clknet_leaf_111_wb_clk_i _02117_ _00785_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13096__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14928_ net1226 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XANTENNA__10303__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10854__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14859_ net1098 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ _04087_ _04089_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09022__X _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16529_ clknet_leaf_82_wb_clk_i _00006_ _01336_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10082__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09001_ _04516_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16693__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13308__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12035__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09527__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ net517 _05419_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11874__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_127_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09834_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\] net754 net702 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__a22o_1
Xfanout558 _07223_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_6
Xfanout569 _07217_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_206_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\] net924 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout562_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ net1061 _04286_ _04316_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__or3b_1
XFILLER_0_69_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09696_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] net778 net732 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a22o_1
XANTENNA__09160__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08647_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net997 vssd1 vssd1 vccd1
+ vccd1 _04276_ sky130_fd_sc_hd__nand2_2
XFILLER_0_178_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout827_A _04512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ _02811_ _04230_ _04227_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08484__A _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10540_ net513 net403 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__nand2_1
XANTENNA__10073__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__X _04400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10471_ _05252_ _05937_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__nand2_1
XANTENNA__10953__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09586__Y _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15110__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04291_ _04292_ _04333_
+ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__nor4_2
X_13190_ team_02_WB.instance_to_wrap.top.pc\[3\] net1024 _02948_ _07337_ vssd1 vssd1
+ vccd1 vccd1 _01484_ sky130_fd_sc_hd__a22o_1
XANTENNA__09766__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net350 net2132 net466 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16797__1341 vssd1 vssd1 vccd1 vccd1 _16797__1341/HI net1341 sky130_fd_sc_hd__conb_1
X_12072_ net354 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\] net471 vssd1
+ vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
Xhold590 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11784__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net408 _06377_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__or2_1
X_15900_ clknet_leaf_16_wb_clk_i _02040_ _00708_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07563__A team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15831_ clknet_leaf_115_wb_clk_i _01971_ _00639_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16720__1352 vssd1 vssd1 vccd1 vccd1 net1352 _16720__1352/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_125_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15762_ clknet_leaf_55_wb_clk_i _01902_ _00570_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12974_ team_02_WB.instance_to_wrap.top.pc\[3\] _05787_ vssd1 vssd1 vccd1 vccd1 _07494_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09151__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14713_ net1097 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
X_11925_ net297 net1960 net484 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
X_15693_ clknet_leaf_49_wb_clk_i _01833_ _00501_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11856_ net310 net1764 net491 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
X_14644_ net1238 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
XFILLER_0_196_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16753__1297 vssd1 vssd1 vccd1 vccd1 _16753__1297/HI net1297 sky130_fd_sc_hd__conb_1
XFILLER_0_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_109_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14575_ net1224 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
X_11787_ net300 net2250 net595 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11261__A1 _04284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16314_ clknet_leaf_51_wb_clk_i _02454_ _01122_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13526_ _03075_ _03086_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__nor2_1
X_10738_ team_02_WB.instance_to_wrap.top.pc\[5\] _06254_ vssd1 vssd1 vccd1 vccd1 _06255_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_70_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13299__X _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11959__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16245_ clknet_leaf_31_wb_clk_i _02385_ _01053_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13457_ _03056_ _03059_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nand2_1
X_10669_ _06128_ _06185_ _04490_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12408_ net641 _07197_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__nand2_8
XFILLER_0_180_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09757__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ net1552 net1013 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[17\]
+ sky130_fd_sc_hd__and2_1
X_16176_ clknet_leaf_23_wb_clk_i _02316_ _00984_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
X_12339_ net362 net2543 net564 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
X_15127_ net1158 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_121_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09509__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_118_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15058_ net1253 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
XFILLER_0_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16096__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ net1098 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
X_07880_ _03581_ _03598_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_182_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09550_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] net868 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13201__A1_N net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ net1048 _04185_ _04194_ _04195_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a31o_1
X_09481_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] net778 net722 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08432_ _04119_ _04131_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08735__C team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ _04060_ _04063_ _04067_ _04070_ _04066_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__a41o_1
XFILLER_0_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10055__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ _03980_ _03990_ _04003_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11869__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout310_A _06840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout408_A _05809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08470__C team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 _06815_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 _06840_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_167_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout777_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 _06955_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_1
Xfanout333 _07013_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_1
XANTENNA__10515__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 _07051_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08479__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net357 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
Xfanout366 _03496_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_2
XANTENNA__09381__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 _06087_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
X_09817_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__inv_2
XANTENNA__09920__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__A3 _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout388 _05901_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_2
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16696__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09748_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\] net751 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] net916 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11710_ net259 net1772 net600 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10294__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15105__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ net298 net2029 net432 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11352__B _06851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ net378 _06567_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14944__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10046__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ net1189 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
X_11572_ net665 net378 _06432_ _07061_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__o31a_1
XANTENNA__09987__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ team_02_WB.instance_to_wrap.top.pc\[4\] net1055 _07064_ net934 vssd1 vssd1
+ vccd1 vccd1 _03005_ sky130_fd_sc_hd__a22o_1
X_10523_ _05782_ net402 vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nor2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_1
XFILLER_0_135_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14291_ net1072 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08178__A1_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16030_ clknet_leaf_4_wb_clk_i _02170_ _00838_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13242_ _06490_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__nor2_1
X_10454_ _04802_ _04822_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input73_A wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08947__B1 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ net976 _07403_ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__or3_1
X_10385_ net547 net385 vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__nor2_1
X_12124_ net284 net1755 net466 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XANTENNA__13299__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ net289 net2119 net470 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
XANTENNA__12403__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ net382 _06513_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__nand2_1
XANTENNA__09372__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09911__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15814_ clknet_leaf_10_wb_clk_i _01954_ _00622_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_16794_ net1338 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__08676__X _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09124__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15745_ clknet_leaf_101_wb_clk_i _01885_ _00553_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12957_ _03294_ _07378_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15015__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10285__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11908_ net243 net1879 net484 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ clknet_leaf_16_wb_clk_i _01816_ _00484_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ net510 _05536_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09013__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14627_ net1134 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
X_16709__1268 vssd1 vssd1 vccd1 vccd1 _16709__1268/HI net1268 sky130_fd_sc_hd__conb_1
X_11839_ net643 _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nand2_4
XFILLER_0_172_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13223__A2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10037__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12431__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11234__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14558_ net1192 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13509_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] _03066_
+ _03067_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__or4_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14489_ net1098 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16228_ clknet_leaf_34_wb_clk_i _02368_ _01036_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16159_ clknet_leaf_62_wb_clk_i _02299_ _00967_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08981_ _04494_ net972 vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__nand2_1
X_07932_ _03613_ _03636_ _03653_ _03654_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12313__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09363__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ _03578_ _03580_ _03583_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__o211a_2
XANTENNA__13492__X _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09602_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\] net922 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a22o_1
X_07794_ _03515_ _03516_ _03513_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_162_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09115__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] net703 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\]
+ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout260_A _06530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10276__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_195_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_195_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ _04113_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_35_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09395_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\] net706 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a22o_1
X_16796__1340 vssd1 vssd1 vccd1 vccd1 _16796__1340/HI net1340 sky130_fd_sc_hd__conb_1
XFILLER_0_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10028__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ _04058_ _03321_ net1007 net2417 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09969__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11599__S net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08277_ _03988_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_78_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout894_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10200__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] net895 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734__1362 vssd1 vssd1 vccd1 vccd1 net1362 _16734__1362/LO sky130_fd_sc_hd__conb_1
Xfanout1106 net1110 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_4
X_16752__1296 vssd1 vssd1 vccd1 vccd1 _16752__1296/HI net1296 sky130_fd_sc_hd__conb_1
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
XANTENNA__12223__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1131 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_4
Xfanout1139 net1141 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_2
XANTENNA__09354__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14939__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13860_ net1149 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11448__A2_N net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ team_02_WB.instance_to_wrap.top.pc\[1\] _04422_ vssd1 vssd1 vccd1 vccd1 _07335_
+ sky130_fd_sc_hd__nand2b_1
X_13791_ net1684 _03278_ net961 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__o21ai_1
X_15530_ clknet_leaf_32_wb_clk_i _01670_ _00338_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12661__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12742_ _06776_ _06797_ net419 vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_210_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12673_ net240 net2014 net432 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15461_ clknet_leaf_28_wb_clk_i _01601_ _00269_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14412_ net1209 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
X_11624_ net379 _07108_ _07110_ net374 _06961_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__o32a_1
XANTENNA__11216__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ clknet_leaf_110_wb_clk_i _01532_ _00200_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11555_ net668 _07031_ _07045_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__o21ai_1
Xwire520 net522 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_2
X_14343_ net1180 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _05124_ _05973_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__nor2_1
X_14274_ net1130 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11486_ _06897_ _06979_ net397 vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13225_ net1470 net1020 net939 _05602_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a22o_1
X_16013_ clknet_leaf_41_wb_clk_i _02153_ _00821_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10437_ _04783_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__or2_1
XANTENNA__12922__A _04489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ _07410_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__xnor2_1
X_10368_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\] _04529_ net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12107_ net2484 net351 net580 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
XANTENNA__12133__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ _07522_ _02862_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__xnor2_1
X_10299_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\] net785 net685 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\]
+ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a221o_1
X_12038_ net354 net2507 net476 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__mux2_1
XANTENNA__14849__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11972__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16777_ net1321 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__09648__A1 _04496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13989_ net1173 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15728_ clknet_leaf_26_wb_clk_i _01868_ _00536_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10258__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15659_ clknet_leaf_15_wb_clk_i _01799_ _00467_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08871__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08200_ _03865_ _03906_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11560__X _07051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09180_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\] net787 net739 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12375__Y _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _03809_ _03817_ _03814_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12308__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10176__X _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08062_ _03758_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__xor2_4
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] net723 _04477_ _04478_
+ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13132__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _03615_ _03618_ _03635_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__a21oi_1
X_08895_ net31 net1029 net986 net2381 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__o22a_1
XANTENNA__14759__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A _07206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _03551_ net329 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_197_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13382__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _03473_ _03496_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__nand2_1
XANTENNA__15501__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11446__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09516_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\] net812 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\]
+ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10249__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\] net725 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08862__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11470__X _06965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A _04524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09378_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\] net815 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08329_ _04035_ _04040_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ net1698 net309 net638 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ _06550_ _06773_ net414 vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__mux2_1
XANTENNA__10961__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13010_ _07455_ _07529_ _07456_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09575__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] net997 _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a22o_1
XANTENNA__11358__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _05625_ _05668_ net551 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16708__1267 vssd1 vssd1 vccd1 vccd1 _16708__1267/HI net1267 sky130_fd_sc_hd__conb_1
XANTENNA__09327__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ net1231 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
X_10084_ _05597_ _05598_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__or3_1
XANTENNA_input36_A gpio_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11792__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\] vssd1 vssd1 vccd1 vccd1
+ net1370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14669__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16700_ net1342 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
X_13912_ net1258 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
XANTENNA__11685__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ net1217 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
XANTENNA__08667__A team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_2
X_16631_ clknet_leaf_95_wb_clk_i _02750_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13843_ net1150 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13426__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16562_ clknet_leaf_90_wb_clk_i _02686_ _01369_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13774_ net1930 _03267_ net960 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__o21ai_1
X_10986_ net1639 net249 net640 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
X_15513_ clknet_leaf_123_wb_clk_i _01653_ _00321_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12725_ _07248_ _07058_ _07031_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16493_ clknet_leaf_81_wb_clk_i _02627_ _01300_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15444_ clknet_leaf_3_wb_clk_i _01584_ _00252_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08606__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ net311 net1767 net435 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ net421 _06750_ _07092_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_170_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12587_ net285 net2328 net438 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__mux2_1
X_15375_ clknet_leaf_84_wb_clk_i _01515_ _00188_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12128__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14326_ net1109 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11538_ net947 _07026_ _07029_ net606 vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__o211a_2
XFILLER_0_111_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11967__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold408 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _06547_ _06853_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__nor2_1
X_14257_ net1222 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_max_cap538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ net633 net938 net1022 net1441 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07746__A team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14188_ net1215 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XANTENNA__09030__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ team_02_WB.instance_to_wrap.top.pc\[12\] net1025 _02906_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01493_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09318__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _03351_ _03386_ _03411_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__and3_1
XFILLER_0_206_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ net1063 _04266_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__nand2_4
XANTENNA_wire610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] _03353_ vssd1 vssd1 vccd1
+ vccd1 _03354_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_179_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11207__S net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 _03302_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09097__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09301_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\] net834 net895 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\]
+ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_192_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09232_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\] net785 net737 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16751__1295 vssd1 vssd1 vccd1 vccd1 _16751__1295/HI net1295 sky130_fd_sc_hd__conb_1
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16733__1361 vssd1 vssd1 vccd1 vccd1 net1361 _16733__1361/LO sky130_fd_sc_hd__conb_1
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09163_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] net807 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ _04679_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08114_ _03795_ _03818_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_211_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_211_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11877__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08045_ _03725_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold920 team_02_WB.instance_to_wrap.top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 net2282
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold931 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13377__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold953 team_02_WB.instance_to_wrap.wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2315
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__B1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__inv_2
XANTENNA__09309__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _04318_ _04339_ _04309_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__a21o_1
XFILLER_0_209_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11667__A1 _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11667__B2 _05356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ net18 net1032 net988 net1696 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ _03532_ _03533_ _03511_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_86_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ net545 net414 vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__or2_2
XANTENNA__09088__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__X _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ net547 net402 vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12510_ net237 net1865 net446 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__mux2_1
X_13490_ team_02_WB.START_ADDR_VAL_REG\[30\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net215 sky130_fd_sc_hd__a21o_1
XFILLER_0_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12441_ net642 _07199_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nand2_2
XFILLER_0_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14952__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12372_ net363 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\] net560 vssd1
+ vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
X_15160_ net1158 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11323_ _05252_ net658 _06113_ _05937_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11787__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14111_ net1108 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
X_15091_ net1111 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09548__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11254_ net837 _06741_ _06751_ net654 _06757_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__o221a_1
X_14042_ net1095 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XANTENNA__11355__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10205_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\] net845 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11185_ _06578_ _06690_ net399 vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\] net754 net734 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__a22o_1
X_16775__1319 vssd1 vssd1 vccd1 vccd1 _16775__1319/HI net1319 sky130_fd_sc_hd__conb_1
X_15993_ clknet_leaf_125_wb_clk_i _02133_ _00801_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07572__Y _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14944_ net1086 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
X_10067_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a22o_1
XANTENNA__12411__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09720__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14875_ net1095 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XANTENNA_clkload1_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16614_ clknet_leaf_87_wb_clk_i _02733_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ net1150 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
XANTENNA__09079__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ clknet_leaf_88_wb_clk_i _02669_ _01352_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09499__Y _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ _03256_ _03257_ _03066_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13280__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ net420 _06481_ _06355_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08826__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15023__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ _06124_ _07231_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16476_ clknet_leaf_70_wb_clk_i net1517 _01284_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
X_13688_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] _03200_ net1642 vssd1 vssd1
+ vccd1 vccd1 _03215_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15427_ clknet_leaf_25_wb_clk_i _01567_ _00235_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12639_ net641 _07210_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09787__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ clknet_leaf_75_wb_clk_i _01498_ _00171_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09251__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14309_ net1114 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
Xhold205 net135 vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 team_02_WB.instance_to_wrap.top.a1.row2\[1\] vssd1 vssd1 vccd1 vccd1 net1578
+ sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ clknet_leaf_70_wb_clk_i _01433_ _00102_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold227 team_02_WB.START_ADDR_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 team_02_WB.instance_to_wrap.top.a1.row1\[9\] vssd1 vssd1 vccd1 vccd1 net1600
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold249 team_02_WB.instance_to_wrap.top.a1.row2\[16\] vssd1 vssd1 vccd1 vccd1 net1611
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11346__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_4
X_09850_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] net817 net887 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\]
+ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a221o_1
Xfanout718 net720 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
Xfanout729 net732 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09691__A _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ net129 net1045 net992 net1375 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
X_09781_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] net755 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a221o_1
XANTENNA__13417__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08732_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__and3_1
XANTENNA__12321__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09711__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__nand2_2
XFILLER_0_178_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07614_ _03326_ _03330_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ net46 net49 net48 net47 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or4b_1
XFILLER_0_163_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13271__B1 _06588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09490__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ _04725_ _04728_ _04730_ _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nor4_2
XFILLER_0_174_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\] net707 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09242__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09077_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] net826 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10805__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1135_X net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ _03744_ _03750_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_96_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15376__Q team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout974_A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11907__Y _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\] net813 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\]
+ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a221o_1
XANTENNA__10540__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ _07481_ _07509_ _07479_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__o21a_1
XANTENNA__08505__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09702__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _04292_ net641 _07201_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__or3_4
XFILLER_0_99_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13851__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14660_ net1132 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
X_11872_ _07190_ _07193_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__nor2_2
XANTENNA__08945__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13611_ _03117_ _03161_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _04928_ net405 vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ net1121 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13262__B1 _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ clknet_leaf_38_wb_clk_i _02470_ _01138_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10076__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13542_ _03078_ _03081_ _03072_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a21oi_1
X_10754_ team_02_WB.instance_to_wrap.top.pc\[29\] _06270_ vssd1 vssd1 vccd1 vccd1
+ _06271_ sky130_fd_sc_hd__and2_1
XANTENNA__09481__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16261_ clknet_leaf_28_wb_clk_i _02401_ _01069_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13473_ team_02_WB.START_ADDR_VAL_REG\[13\] net1071 net1005 vssd1 vssd1 vccd1 vccd1
+ net196 sky130_fd_sc_hd__a21o_1
X_10685_ team_02_WB.instance_to_wrap.top.pc\[13\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _06202_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15212_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[3\]
+ _00025_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09769__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ net303 net2533 net457 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__mux2_1
XANTENNA__09776__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16192_ clknet_leaf_18_wb_clk_i _02332_ _01000_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15143_ net1156 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XANTENNA__11040__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net272 net2346 net562 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__mux2_1
XANTENNA__12406__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13317__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _06195_ _06212_ _06213_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__nand3_1
X_12286_ net282 net2150 net571 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__mux2_1
X_15074_ net1245 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
X_14025_ net1216 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
X_11237_ _05127_ _05943_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10000__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ _04996_ net664 _06667_ net795 _06668_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__o221a_1
X_16732__1360 vssd1 vssd1 vccd1 vccd1 net1360 _16732__1360/LO sky130_fd_sc_hd__conb_1
X_16750__1294 vssd1 vssd1 vccd1 vccd1 _16750__1294/HI net1294 sky130_fd_sc_hd__conb_1
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\] net813 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ _05630_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a221o_1
XANTENNA__12141__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10450__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ net415 _06107_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__or2_1
X_15976_ clknet_leaf_25_wb_clk_i _02116_ _00784_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14927_ net1199 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11980__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14858_ net1179 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XANTENNA__10854__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13480__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ net1154 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ net1114 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10067__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16528_ clknet_leaf_82_wb_clk_i _00005_ _01335_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16459_ clknet_leaf_84_wb_clk_i net1570 _01267_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
X_09000_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ _04499_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09224__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_wb_clk_i_X clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10625__A team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09902_ net971 net624 net544 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12840__A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09932__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09833_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\] net786 net718 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__a221o_1
Xfanout559 _07223_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_4
XANTENNA_fanout290_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Right_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_206_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08999__C_N net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12051__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10360__A _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\] net806 net880 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__a221o_1
X_08715_ _04338_ _04340_ _04341_ _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__and4b_1
X_09695_ _05207_ _05209_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nor2_1
XANTENNA__11890__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08646_ _04265_ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ net1637 _04240_ _04225_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout722_A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_X net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09999__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16774__1318 vssd1 vssd1 vccd1 vccd1 _16774__1318/HI net1318 sky130_fd_sc_hd__conb_1
XFILLER_0_45_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470_ _05231_ _05251_ _05291_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a21o_1
XANTENNA__08635__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\] net906 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ _04645_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a221o_1
XANTENNA__12226__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ net362 net2154 net466 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10230__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08005__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ net360 net2274 net472 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
Xhold580 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _06531_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__xnor2_1
X_15830_ clknet_leaf_22_wb_clk_i _01970_ _00638_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_204_Left_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15761_ clknet_leaf_0_wb_clk_i _01901_ _00569_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12973_ team_02_WB.instance_to_wrap.top.pc\[3\] _05787_ vssd1 vssd1 vccd1 vccd1 _07493_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10297__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14712_ net1195 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
X_11924_ net310 net1961 net483 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
X_15692_ clknet_leaf_2_wb_clk_i _01832_ _00500_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14643_ net1073 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
X_11855_ net300 net1774 net493 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10049__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _06320_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14574_ net1073 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
XFILLER_0_200_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11786_ net294 net2072 net594 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16313_ clknet_leaf_125_wb_clk_i _02453_ _01121_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10737_ team_02_WB.instance_to_wrap.top.pc\[4\] team_02_WB.instance_to_wrap.top.pc\[3\]
+ team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16244_ clknet_leaf_3_wb_clk_i _02384_ _01052_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15885__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13456_ _03038_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__or2_1
XANTENNA__08653__B_N team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10668_ net995 _05580_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_1
XANTENNA__09206__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12407_ net348 net1919 net458 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16175_ clknet_leaf_42_wb_clk_i _02315_ _00983_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12136__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10599_ _04462_ _06114_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__or2_4
X_13387_ net2477 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[16\]
+ sky130_fd_sc_hd__and2_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126_ net1165 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
X_12338_ net355 net2421 net566 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15057_ net1254 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
X_12269_ net340 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net575 vssd1
+ vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09914__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ net1195 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_182_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09017__Y _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15265__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ clknet_leaf_120_wb_clk_i _02099_ _00767_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14587__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ team_02_WB.instance_to_wrap.top.a1.row1\[17\] _04186_ vssd1 vssd1 vccd1 vccd1
+ _04195_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09480_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_201_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08431_ _04119_ _04131_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13226__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _04060_ _04063_ _04070_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and3_1
XFILLER_0_191_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09445__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11252__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08293_ _03948_ _03967_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12835__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10626__Y _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12046__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11738__X _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _06815_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_1
XFILLER_0_10_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 net315 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_2
Xfanout323 _06955_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout334 _06994_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XANTENNA_fanout672_A _04469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10515__B2 _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _07051_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_1
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
X_09816_ net970 net626 net543 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__o21ai_1
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_2
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout389 net392 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_2
X_09747_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\] net844 _05261_ _05262_
+ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13465__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_190_Right_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] net819 net904 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__a221o_1
XANTENNA__09684__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08629_ net97 net1521 net955 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XANTENNA__11491__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13323__A1_N team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11640_ net2039 net353 net637 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09436__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _05738_ _06110_ net657 _05737_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_64_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ net1439 net983 net965 _03004_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__a22o_1
X_10522_ net498 net402 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14290_ net1184 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08661__C _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10453_ _04802_ _04822_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and2_1
X_13241_ _06523_ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10265__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08947__A1 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ net403 vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__inv_2
XANTENNA_input66_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ _07387_ _07401_ _07402_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__and3_1
XANTENNA__11795__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ net275 net2347 net467 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
X_12054_ net276 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\] net470 vssd1
+ vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
X_11005_ net420 _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input21_X net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net893 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_8
X_15813_ clknet_leaf_28_wb_clk_i _01953_ _00621_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_16793_ net1337 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
X_15744_ clknet_leaf_18_wb_clk_i _01884_ _00552_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12956_ _03294_ _07378_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__nand2_1
XANTENNA__09675__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11907_ _04452_ _07199_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__nand2_4
X_15675_ clknet_leaf_34_wb_clk_i _01815_ _00483_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _07404_ _07406_ _07386_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_47_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14626_ net1129 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
X_11838_ _07188_ _07193_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09427__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14557_ net1181 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XANTENNA__09948__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ net353 net2270 net596 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__mux2_1
XANTENNA__10727__X _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\]
+ _03065_ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14488_ net1197 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16227_ clknet_leaf_26_wb_clk_i _02367_ _01035_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13439_ _03043_ _03044_ _03040_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08938__A1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ clknet_leaf_5_wb_clk_i _02298_ _00966_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09060__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15109_ net1102 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16089_ clknet_leaf_123_wb_clk_i _02229_ _00897_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_08980_ _04491_ _04493_ net972 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__and3_4
X_07931_ _03575_ _03612_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07862_ _03549_ _03572_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_208_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09601_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] net805 _05104_ _05117_
+ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a211o_1
X_16773__1317 vssd1 vssd1 vccd1 vccd1 _16773__1317/HI net1317 sky130_fd_sc_hd__conb_1
X_07793_ _03451_ _03478_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_162_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] net755 net747 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09666__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _04973_ _04975_ _04979_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout253_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08414_ _04119_ _04120_ _04115_ _04116_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09394_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] net743 net724 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13137__A2_N net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09418__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08345_ _04050_ _04051_ _04057_ _04043_ _04037_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_46_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08276_ _03962_ _03987_ _03964_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1270_A team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_X net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1107 net1110 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1129 net1131 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_111_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_199_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _04422_ team_02_WB.instance_to_wrap.top.pc\[1\] vssd1 vssd1 vccd1 vccd1 _07334_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_202_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13790_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] _03278_
+ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__and2_1
XANTENNA__14020__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09657__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08656__C _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ net380 _06550_ _07001_ _07262_ _07264_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__o2111a_1
XANTENNA__14955__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15460_ clknet_leaf_36_wb_clk_i _01600_ _00268_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12672_ net641 _07212_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__nand2_8
XANTENNA__09409__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14411_ net1125 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
X_11623_ net390 _06039_ _06042_ _07109_ net395 vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__o311a_1
X_15391_ clknet_leaf_61_wb_clk_i _01531_ _00199_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08672__B team_02_WB.instance_to_wrap.top.a1.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14342_ net1204 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
X_11554_ net836 _07032_ _07039_ _06117_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_146_Left_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire532 _05102_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09290__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10975__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10505_ _04994_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14273_ net1258 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
X_11485_ _06938_ _06978_ net367 vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold887_X net2249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16012_ clknet_leaf_126_wb_clk_i _02152_ _00820_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13224_ net1475 net1022 net939 _05555_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__a22o_1
X_10436_ _05950_ _05952_ _04823_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12922__B _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ _07384_ _07385_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__or2_1
X_10367_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] net922 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a22o_1
XANTENNA__12414__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12106_ net1679 net364 net580 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
X_10298_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\] net757 net741 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__a22o_1
X_13086_ _07461_ _07462_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13141__A2 _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ net360 net2169 net477 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_155_Left_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09896__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16776_ net1320 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
X_13988_ net1098 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XANTENNA__09648__A2 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ clknet_leaf_41_wb_clk_i _01867_ _00535_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12939_ team_02_WB.instance_to_wrap.top.pc\[22\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _07459_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15658_ clknet_leaf_37_wb_clk_i _01798_ _00466_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ net1229 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_164_Left_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15589_ clknet_leaf_29_wb_clk_i _01729_ _00397_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ _03809_ _03814_ _03817_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09281__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09820__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08061_ _03709_ _03740_ _03710_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11288__X _06791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12324__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10194__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\] net782 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_173_Left_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07914_ _03632_ _03634_ _03621_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a21o_1
XANTENNA__13944__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ net32 net1032 net988 team_02_WB.instance_to_wrap.ramload\[8\] vssd1 vssd1
+ vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XANTENNA__09887__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ _03558_ _03566_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout370_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07776_ _03465_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_88_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09515_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] net923 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\] net761 net677 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_182_Left_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09377_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\] net877 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout802_A _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10808__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08492__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08328_ _04030_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09272__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15379__Q team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _03925_ _03960_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _06664_ _06772_ net399 vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10221_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and2b_2
XFILLER_0_30_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12234__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] net649 _05668_ vssd1
+ vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a21o_1
XANTENNA__11358__B _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14960_ net1227 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
X_10083_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\] net857 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a221o_1
XANTENNA__12331__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\] vssd1 vssd1 vccd1 vccd1
+ net1371 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ net1233 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XANTENNA__11685__A2 _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ net1124 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ clknet_leaf_95_wb_clk_i _02749_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10893__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ net1150 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16561_ clknet_leaf_90_wb_clk_i _02685_ _01368_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08838__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\]
+ _03265_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__and3_1
XANTENNA__11437__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ net604 _06491_ _06497_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__and3_2
XFILLER_0_186_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15512_ clknet_leaf_122_wb_clk_i _01652_ _00320_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12724_ _05833_ net668 _07075_ _07175_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16492_ clknet_leaf_92_wb_clk_i _02626_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08683__A team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15443_ clknet_leaf_52_wb_clk_i _01583_ _00251_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12655_ net302 net2560 net437 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12409__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11606_ net421 _06749_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__nor2_1
X_15374_ clknet_leaf_85_wb_clk_i _01514_ _00187_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_12586_ net273 net2535 net441 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__mux2_1
XANTENNA__09802__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10948__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14325_ net1257 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16772__1316 vssd1 vssd1 vccd1 vccd1 _16772__1316/HI net1316 sky130_fd_sc_hd__conb_1
X_11537_ team_02_WB.instance_to_wrap.top.pc\[6\] net974 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\]
+ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12933__A team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_150_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ net1232 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
X_11468_ net376 _06773_ _06961_ net383 _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__a221o_1
XANTENNA__08622__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ _04821_ net936 net1020 net1388 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a2bb2o_1
X_10419_ net610 _05251_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nor2_1
XANTENNA__10453__A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14187_ net1098 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XANTENNA__11373__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _06847_ _06896_ net369 vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13138_ _04280_ _02904_ _02905_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11983__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13069_ _07430_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__xnor2_1
Xhold1109 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09869__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13169__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03349_ vssd1 vssd1 vccd1
+ vccd1 _03353_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_179_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07561_ net1 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__inv_2
XANTENNA__08829__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16759_ net1303 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
X_09300_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\] net811 net891 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10100__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09231_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\] net757 net729 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12319__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09162_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\] net904 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09254__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08113_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13107__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09093_ _04588_ _04608_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_211_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12843__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08044_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03722_ vssd1 vssd1 vccd1
+ vccd1 _03766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold910 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold921 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold932 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12054__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold965 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1125_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _05489_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout585_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08946_ _04318_ _04339_ _04309_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11116__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__A2 _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ net19 net1031 _04432_ net1590 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout752_A _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07828_ _03546_ _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_190_Left_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07759_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ net498 net385 _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09493__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ _04934_ _04941_ _04944_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__or4_4
XANTENNA__12229__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ net349 net2121 net454 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__mux2_1
XANTENNA__09245__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ net355 net2375 net561 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ net1188 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
X_11322_ _06821_ _06822_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__nor2_1
X_15090_ net1072 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14041_ net1089 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
X_11253_ _05127_ net663 _06754_ net795 _06755_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__o221a_1
XANTENNA__10158__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__B2 _06854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\] net747 net692 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__a22o_1
X_11184_ _06629_ _06689_ net371 vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10135_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\] net691 _05650_ _05651_
+ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a211o_1
XFILLER_0_207_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15992_ clknet_leaf_120_wb_clk_i _02132_ _00800_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11107__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14943_ net1109 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
X_10066_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14874_ net1096 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08965__X _04482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10330__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16613_ clknet_leaf_92_wb_clk_i _02732_ _01406_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13825_ net1149 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16544_ clknet_leaf_87_wb_clk_i _02668_ _01351_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13756_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o211a_1
X_10968_ net410 _06480_ _06359_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__o21a_1
XANTENNA__08617__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09484__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ _04355_ _06163_ _06249_ _07123_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__o22a_1
X_16475_ clknet_leaf_69_wb_clk_i net1483 _01283_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13687_ net1592 _03200_ _03214_ net1141 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12139__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10899_ _06413_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__inv_2
XFILLER_0_183_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15426_ clknet_leaf_115_wb_clk_i _01566_ _00234_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12638_ net2085 net347 net552 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09236__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11978__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ clknet_leaf_75_wb_clk_i _01497_ _00170_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12569_ net356 net2276 net445 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14308_ net1137 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15288_ clknet_leaf_72_wb_clk_i _01432_ _00101_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold206 _02601_ vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 team_02_WB.START_ADDR_VAL_REG\[31\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 team_02_WB.instance_to_wrap.ramload\[25\] vssd1 vssd1 vccd1 vccd1 net1590
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold239 team_02_WB.instance_to_wrap.ramload\[1\] vssd1 vssd1 vccd1 vccd1 net1601
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ net1115 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13197__C _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10149__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09972__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout708 _04387_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_4
Xfanout719 net720 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
X_08800_ net1427 net1045 net991 team_02_WB.instance_to_wrap.ramaddr\[31\] vssd1 vssd1
+ vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
X_09780_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] net772 net696 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a22o_1
XANTENNA__12602__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08731_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08662_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__nand2_2
XANTENNA__10321__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07613_ _03332_ _03335_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ net52 net51 net54 net53 vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__or4_1
XANTENNA__13031__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09475__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13271__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12049__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout333_A _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] net891 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\]
+ _04716_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09227__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13023__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11888__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09145_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\] net788 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1242_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09076_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] net900 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\]
+ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11189__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ _03712_ _03738_ _03749_ _03745_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_96_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold740 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold751 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1128_X net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold773 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09978_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\] net867 net857 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a22o_1
XANTENNA__12512__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] net1009 _04447_ _04448_ vssd1
+ vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11940_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] _04333_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or3b_4
XFILLER_0_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16771__1315 vssd1 vssd1 vccd1 vccd1 _16771__1315/HI net1315 sky130_fd_sc_hd__conb_1
XFILLER_0_207_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11871_ net348 net2303 net490 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _03289_ net1049 _03127_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__nor3_1
XANTENNA__11652__A _04482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10822_ _04971_ net388 vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ net1189 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13262__A1 _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09466__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ _03078_ _03086_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__nor2_1
X_10753_ team_02_WB.instance_to_wrap.top.pc\[28\] team_02_WB.instance_to_wrap.top.pc\[27\]
+ _06269_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__and3_1
X_16260_ clknet_leaf_32_wb_clk_i _02400_ _01068_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input96_A wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ team_02_WB.START_ADDR_VAL_REG\[12\] net1070 net1004 vssd1 vssd1 vccd1 vccd1
+ net195 sky130_fd_sc_hd__a21o_1
X_10684_ team_02_WB.instance_to_wrap.top.pc\[13\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _06201_ sky130_fd_sc_hd__nand2_1
X_15211_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[2\]
+ _00024_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11798__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ net292 net2341 net455 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16191_ clknet_leaf_60_wb_clk_i _02331_ _00999_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10379__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15142_ net1156 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12354_ net288 net2152 net560 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XANTENNA__11099__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _06800_ _06803_ _06806_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_39_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13317__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15073_ net1168 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12285_ net269 net2497 net570 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__mux2_1
XANTENNA__11328__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ net1113 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
X_11236_ net1648 net272 net639 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12930__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net423 _06673_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__nand2_1
XANTENNA__12422__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\] net817 net907 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\]
+ _05631_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__a221o_1
X_15975_ clknet_leaf_38_wb_clk_i _02115_ _00783_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11098_ net411 _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14926_ net1083 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
X_10049_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] net717 net838 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10303__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14857_ net1210 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ net1142 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14788_ net1136 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XANTENNA__09457__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ _03245_ _03246_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16527_ clknet_leaf_84_wb_clk_i _02660_ _01334_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.busy_o
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09209__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16458_ clknet_leaf_43_wb_clk_i net1401 _01266_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15409_ clknet_leaf_128_wb_clk_i _01549_ _00217_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_154_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16389_ clknet_leaf_89_wb_clk_i _02524_ _01197_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11501__S net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13308__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09901_ _05405_ _05412_ _05415_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nor4_2
XFILLER_0_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13428__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] net710 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12332__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] net830 net887 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout283_A _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _04311_ _04276_ _04320_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__mux2_1
XANTENNA__13952__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09694_ _05207_ _05209_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__or2_1
XANTENNA__09696__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09160__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08645_ _04271_ _04273_ _04268_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout450_A _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09448__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ _04180_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__nor2_1
XANTENNA__10359__Y _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13399__A team_02_WB.instance_to_wrap.ramload\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] net890 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\] net735 net844 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12070_ net345 net2153 net471 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
Xhold570 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 team_02_WB.instance_to_wrap.ramload\[26\] vssd1 vssd1 vccd1 vccd1 net1943
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _04863_ _05950_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__nor2_1
XANTENNA__13180__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ clknet_leaf_23_wb_clk_i _01900_ _00568_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12972_ _07490_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__and2_1
XANTENNA__09687__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1 net2632
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net300 net2348 net485 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__mux2_1
XANTENNA__09151__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ net1208 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15691_ clknet_leaf_15_wb_clk_i _01831_ _00499_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14642_ net1184 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XANTENNA__09439__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13235__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ net295 net1868 net492 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10805_ _04842_ net405 vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14573_ net1128 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
X_11785_ net284 net1816 net592 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16312_ clknet_leaf_122_wb_clk_i _02452_ _01120_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13524_ _03073_ _03077_ _03061_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ _06245_ net652 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] net496
+ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12925__B _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16243_ clknet_leaf_56_wb_clk_i _02383_ _01051_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ _03036_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__nand2_1
XANTENNA__12417__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ _06128_ _06183_ _04490_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a21oi_4
X_12406_ net351 net1920 net458 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
X_16174_ clknet_leaf_46_wb_clk_i _02314_ _00982_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13386_ team_02_WB.instance_to_wrap.ramload\[15\] net1014 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[15\] sky130_fd_sc_hd__and2_1
XANTENNA__09611__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ _04462_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__nor2_1
X_15125_ net1163 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
X_12337_ net358 net2120 net565 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_50_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15056_ net1263 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XANTENNA__08630__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ net333 net1720 net575 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14007_ net1207 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15029__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ _05081_ _06113_ _06116_ _05082_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__o22a_1
XANTENNA__12152__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net322 net2227 net576 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11991__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09678__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15958_ clknet_leaf_22_wb_clk_i _02098_ _00766_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09142__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ net1204 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
X_15889_ clknet_leaf_0_wb_clk_i _02029_ _00697_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09033__Y _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ _04042_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08292_ _03969_ _04002_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09850__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12835__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13529__A2 _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12327__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14108__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09602__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16770__1314 vssd1 vssd1 vccd1 vccd1 _16770__1314/HI net1314 sky130_fd_sc_hd__conb_1
XFILLER_0_42_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13947__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12851__A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12062__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout313 net315 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout324 _06955_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout335 _06994_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1205_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_2
X_09815_ _05325_ _05328_ _05329_ _05331_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__nor4_1
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 _07087_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09381__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 net373 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_2
Xfanout379 net381 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_2
XFILLER_0_185_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] net767 net703 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\]
+ _05253_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__a221o_1
XANTENNA__13465__A1 team_02_WB.START_ADDR_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\] net888 net868 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout832_A _04506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ net98 team_02_WB.START_ADDR_VAL_REG\[4\] net957 vssd1 vssd1 vccd1 vccd1 _02632_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08892__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04169_ vssd1 vssd1 vccd1
+ vccd1 _04228_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_59_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11570_ _05736_ net660 net654 _07056_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09841__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10521_ _04461_ _05963_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08942__C _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12237__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ _06556_ _06588_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__nand2b_1
X_10452_ _04713_ _04733_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__A2 _04339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07604__C1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13171_ net229 _07502_ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__nand3_1
X_10383_ _04422_ net968 _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12122_ net288 net1929 net469 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XANTENNA_input59_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12053_ net282 net2127 net471 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__mux2_1
X_11004_ _06514_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__and2_1
XANTENNA__09372__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__X _07150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 _04538_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_8
X_15812_ clknet_leaf_34_wb_clk_i _01952_ _00620_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout891 net893 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12700__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ net1336 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__08686__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15743_ clknet_leaf_58_wb_clk_i _01883_ _00551_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12955_ _07473_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _06280_ _07193_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15674_ clknet_leaf_52_wb_clk_i _01814_ _00482_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12886_ _07386_ _07405_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11219__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14625_ net1260 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
X_11837_ net346 net2571 net588 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ net1191 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
X_11768_ net364 net1842 net596 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__mux2_1
XANTENNA__08625__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09832__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ _03064_ _03068_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10719_ team_02_WB.instance_to_wrap.top.pc\[26\] _06147_ _06235_ vssd1 vssd1 vccd1
+ vccd1 _06236_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16208__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14487_ net1210 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ net1001 net995 _07123_ team_02_WB.instance_to_wrap.top.pc\[0\] vssd1 vssd1
+ vccd1 vccd1 _07185_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_151_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13438_ _03043_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__nand2_1
X_16226_ clknet_leaf_119_wb_clk_i _02366_ _01034_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11986__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08938__A2 _04346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ clknet_leaf_10_wb_clk_i _02297_ _00965_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13369_ net1623 team_02_WB.instance_to_wrap.top.ru.next_iready vssd1 vssd1 vccd1
+ vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[31\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_184_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15108_ net1072 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
X_16088_ clknet_leaf_114_wb_clk_i _02228_ _00896_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_07930_ _03612_ _03613_ _03636_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a21oi_2
X_15039_ net1244 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XANTENNA__09899__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14598__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\] net828 net905 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\]
+ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12610__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07792_ _03490_ _03491_ _03492_ net366 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09531_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\] net724 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09115__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11458__B1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] net816 _04976_ _04978_
+ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a211o_1
XFILLER_0_188_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08874__B2 team_02_WB.instance_to_wrap.ramload\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_148_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08413_ _04119_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_195_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09393_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] net767 net759 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12846__A _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08344_ _04040_ _04052_ _04024_ _04035_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__and4b_1
XFILLER_0_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09823__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08275_ net2478 net1007 net980 _03990_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
XANTENNA__12057__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1155_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11896__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1110 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1171 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09354__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12520__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11449__B1 _06943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\] net829 net879 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\]
+ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ net380 _06347_ _06407_ _06453_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08656__D net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10121__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ net348 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\] net434 vssd1
+ vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10828__X _06344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14410_ net1176 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
X_11622_ net389 _07071_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__nand2_1
XANTENNA__08617__A1 team_02_WB.START_ADDR_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15390_ clknet_leaf_5_wb_clk_i _01530_ _00198_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09814__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ net1113 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
X_11553_ net794 _07040_ _07041_ net665 _07043_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10975__A2 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire533 _04841_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_42_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504_ _04970_ _04992_ _05039_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__o21ai_1
X_14272_ net1102 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
X_11484_ _06298_ _06300_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
X_16011_ clknet_leaf_15_wb_clk_i _02151_ _00819_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13223_ net1537 _00012_ net939 _05510_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10435_ _04863_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__or2_1
XANTENNA__10188__B1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09593__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ net229 _07507_ _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10366_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] net926 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a22o_1
X_12105_ net2515 net354 net582 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
X_13085_ net1027 _02861_ net1025 team_02_WB.instance_to_wrap.top.pc\[21\] vssd1 vssd1
+ vccd1 vccd1 _01502_ sky130_fd_sc_hd__a2bb2o_1
X_10297_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\] net689 net842 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a22o_1
X_12036_ net343 net2329 net476 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12430__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16775_ net1319 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
X_13987_ net1137 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15726_ clknet_leaf_47_wb_clk_i _01866_ _00534_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10112__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ team_02_WB.instance_to_wrap.top.pc\[22\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _07458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15657_ clknet_leaf_112_wb_clk_i _01797_ _00465_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12869_ _05788_ net498 vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_177_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14608_ net1232 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15588_ clknet_leaf_35_wb_clk_i _01728_ _00396_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09805__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14539_ net1124 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14881__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_190_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ _03771_ _03776_ _03781_ _03759_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12672__Y _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16209_ clknet_leaf_0_wb_clk_i _02349_ _01017_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10179__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12605__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09584__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08962_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\] net727 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_164_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07913_ _03632_ _03634_ _03621_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a21oi_2
X_08893_ net33 net1029 net986 net2230 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12340__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ _03530_ _03559_ _03532_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_197_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07775_ _03474_ net366 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout363_A _07107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09514_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] net907 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09445_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] net737 _04952_ _04955_
+ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\] net925 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08327_ _04038_ _04031_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11603__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08258_ _03910_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12515__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ _03876_ _03896_ _03867_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10220_ net422 net502 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13200__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09575__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] _04330_ vssd1 vssd1
+ vccd1 vccd1 _05668_ sky130_fd_sc_hd__and2_1
XANTENNA__08788__X _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10082_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\] net910 net890 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a22o_1
X_13910_ net1258 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12250__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ net1179 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
X_13841_ net1150 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13772_ _03267_ _03268_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__nor2_1
X_16560_ clknet_leaf_87_wb_clk_i _02684_ _01367_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ net974 _06493_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__a21o_1
X_15511_ clknet_leaf_122_wb_clk_i _01651_ _00319_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12723_ _06283_ _07246_ _06375_ _05961_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_44_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16491_ clknet_leaf_80_wb_clk_i net1057 _01299_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08683__B team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12654_ net293 net1793 net435 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__mux2_1
X_15442_ clknet_leaf_54_wb_clk_i _01582_ _00250_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11605_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12585_ net288 net2038 net438 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__mux2_1
X_15373_ clknet_leaf_85_wb_clk_i _01513_ _00186_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10948__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input81_X net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14324_ net1239 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
X_11536_ net1000 _07027_ net947 vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12933__B _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ net1220 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
X_11467_ net413 _06549_ net424 vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12425__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13206_ _04774_ net936 net1020 net1407 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10418_ _05294_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08470__A_N team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14186_ net1118 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
X_11398_ _06305_ _06307_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13137_ _06911_ net234 net231 _02903_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__a2bb2o_1
X_10349_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] net705 net701 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09318__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ _07361_ _07362_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__and2b_1
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ net280 net1916 net477 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XANTENNA__12160__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10333__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire429_A _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07560_ net1140 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__inv_2
X_16758_ net1302 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_158_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ clknet_leaf_13_wb_clk_i _01849_ _00517_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16689_ clknet_leaf_71_wb_clk_i _02806_ _01413_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09230_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\] net725 _04736_ _04739_
+ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_118_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10628__B _06143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09161_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\] net885 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\]
+ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08112_ _03792_ _03830_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09092_ _04588_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_211_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08043_ _03763_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__and2_1
Xhold900 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12335__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold911 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09557__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10363__B _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold955 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11364__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold977 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13955__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1020_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _05491_ _05510_ net968 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__mux2_2
Xhold999 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1118_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _04458_ _04460_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_110_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout578_A _07214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ net20 net1032 net988 net1943 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XANTENNA__10324__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _03549_ _03547_ _03536_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__and3b_1
XANTENNA__14786__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ _03416_ _03479_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07689_ _03393_ _03394_ _03377_ _03384_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout912_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15913__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09428_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\] net915 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\]
+ _04932_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09359_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] net768 _04874_ _04875_
+ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13214__A1_N net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12370_ net358 net2047 net562 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11321_ net411 _06107_ net419 vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_185_Right_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12245__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ net1196 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
XANTENNA__09548__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ _05123_ net662 _06753_ _06037_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__a22o_1
XANTENNA__08024__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\] net724 _05718_ _05719_
+ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a211o_1
XANTENNA__16419__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11183_ _06688_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__inv_2
XANTENNA_input41_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] net775 net763 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a22o_1
X_15991_ clknet_leaf_120_wb_clk_i _02131_ _00799_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11107__A2 _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11385__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14942_ net1128 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
X_10065_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net791 net650 _05581_
+ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_128_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09181__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09720__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14873_ net1088 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16612_ clknet_leaf_91_wb_clk_i _02731_ _01405_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_199_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ net1147 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16543_ clknet_leaf_82_wb_clk_i _00015_ _01350_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10967_ net407 _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__or2_1
X_13755_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\] vssd1 vssd1 vccd1
+ vccd1 _03256_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13280__A2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11291__A1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ net72 team_02_WB.EN_VAL_REG _07230_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__mux2_1
XANTENNA__10094__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16474_ clknet_leaf_69_wb_clk_i net1485 _01282_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
X_10898_ _06032_ _06373_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__xor2_1
X_13686_ _03200_ _03204_ net1592 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_174_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09796__Y _05313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15425_ clknet_leaf_102_wb_clk_i _01565_ _00233_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12637_ net1657 net352 net552 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11579__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09787__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ net359 net2604 net444 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__mux2_1
X_15356_ clknet_leaf_74_wb_clk_i _01496_ _00169_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_156_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ net1137 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
X_11519_ net953 _07010_ _07011_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__or3_1
XANTENNA__12155__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10464__A _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ net331 net2131 net557 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__mux2_1
X_15287_ clknet_leaf_82_wb_clk_i _01431_ _00100_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold207 net106 vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_02_WB.instance_to_wrap.top.a1.row2\[0\] vssd1 vssd1 vccd1 vccd1 net1580
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold229 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ net1190 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XANTENNA__13197__D _04289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11346__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ net1087 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
Xfanout709 net712 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08730_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] net931 vssd1 vssd1 vccd1
+ vccd1 _04359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10306__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09172__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ net1060 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] _04286_ vssd1
+ vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__or3_1
XANTENNA__09711__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03331_ _03333_ vssd1 vssd1
+ vccd1 vccd1 _03335_ sky130_fd_sc_hd__or3_1
X_08592_ net50 net39 net64 _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12838__B _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10198__X _05715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09475__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13271__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] net928 net811 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12854__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13023__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout326_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09144_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\] net844 _04654_ _04658_
+ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1068_A _00018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] net908 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12065__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ _03720_ _03728_ _03731_ _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_112_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold730 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold741 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout695_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold752 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 team_02_WB.instance_to_wrap.top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 net2125
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold785 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 team_02_WB.instance_to_wrap.ramload\[20\] vssd1 vssd1 vccd1 vccd1 net2158
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\] net833 net804 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\]
+ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout862_A _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net1047 _04218_ _04232_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09163__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10848__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10848__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ net166 net1043 net1035 net1394 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ net352 net1776 net490 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821_ _05017_ net404 _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11652__B _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10076__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13540_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] _03061_ _03097_ _03098_
+ net1068 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__o221a_1
X_10752_ team_02_WB.instance_to_wrap.top.pc\[26\] _06268_ vssd1 vssd1 vccd1 vccd1
+ _06269_ sky130_fd_sc_hd__and2_1
X_13471_ team_02_WB.START_ADDR_VAL_REG\[11\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net194 sky130_fd_sc_hd__a21o_1
XFILLER_0_180_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10683_ net789 _05785_ _06127_ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__o22a_2
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12422_ net286 net1700 net455 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
X_15210_ clknet_leaf_88_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[1\]
+ _00023_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09769__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16190_ clknet_leaf_1_wb_clk_i _02330_ _00998_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input89_A wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ net279 net1771 net560 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
X_15141_ net1142 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11304_ net670 _06792_ _06805_ net837 vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__o2bb2a_1
X_15072_ net1166 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
X_12284_ net261 net2378 net570 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14023_ net1181 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11235_ net606 _06732_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__and3_4
XANTENNA__12703__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _06401_ _06665_ net413 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10290__Y _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] net882 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__a22o_1
X_11097_ _06479_ _06605_ net399 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__mux2_1
X_15974_ clknet_leaf_6_wb_clk_i _02114_ _00782_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10048_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\] net677 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a22o_1
X_14925_ net1126 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12939__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold90 _02566_ vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
X_14856_ net1117 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XANTENNA__08628__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ net1162 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14787_ net1134 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
X_11999_ net334 net2147 net480 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XANTENNA__11054__S net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16526_ clknet_leaf_1_wb_clk_i _00016_ _01333_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dfrtp_2
XANTENNA__10067__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ net2563 _03244_ net950 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11989__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16457_ clknet_leaf_44_wb_clk_i net1387 _01265_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13669_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_116_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11016__A1 _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15408_ clknet_leaf_30_wb_clk_i _01548_ _00216_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_154_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13489__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11016__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16388_ clknet_leaf_89_wb_clk_i _02523_ _01196_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15339_ clknet_leaf_42_wb_clk_i _01482_ _00152_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09900_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] net914 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\]
+ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a221o_1
XANTENNA__12613__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] net751 _05338_ _05341_
+ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_169_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\] net814 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_206_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09145__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__inv_2
X_09693_ net523 _05206_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08644_ net1061 _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08575_ team_02_WB.instance_to_wrap.top.a1.hexop\[4\] _04231_ _04228_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_25_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout443_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10058__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11899__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09127_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] net820 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\]
+ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a221o_1
XANTENNA__08959__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09058_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] net751 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a22o_1
XANTENNA__10230__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ _03726_ _03727_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12523__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold571 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _05970_ _05971_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09384__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16499__Q team_02_WB.START_ADDR_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ team_02_WB.instance_to_wrap.top.pc\[4\] _05742_ vssd1 vssd1 vccd1 vccd1 _07491_
+ sky130_fd_sc_hd__or2_1
Xhold1260 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net2633
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ net1084 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
XANTENNA__10297__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ net292 net2164 net483 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__mux2_1
X_15690_ clknet_leaf_39_wb_clk_i _01830_ _00498_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14641_ net1222 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
X_11853_ net285 net1853 net490 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10049__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ _04886_ net388 vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14572_ net1215 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XFILLER_0_200_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11784_ net274 net2598 net595 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08972__A _04482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16311_ clknet_leaf_115_wb_clk_i _02451_ _01119_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ _03077_ _03081_ _03083_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_171_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ _06161_ _06251_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16242_ clknet_leaf_18_wb_clk_i _02382_ _01050_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13454_ _03032_ _02763_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__or2_1
X_10666_ net994 _05441_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12405_ net364 net2325 net458 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__mux2_1
X_16173_ clknet_leaf_49_wb_clk_i _02313_ _00981_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13385_ net1533 net1013 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[14\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10597_ _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__or2_2
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15124_ net1165 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
X_12336_ net343 net2578 net566 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
XANTENNA__08911__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12267_ net334 net1719 net574 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12433__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15055_ net1250 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XANTENNA__09375__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__inv_2
X_14006_ net1106 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XANTENNA__09914__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12198_ net317 net2380 net576 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11149_ net605 _06649_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_182_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09127__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ clknet_leaf_22_wb_clk_i _02097_ _00765_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15045__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10288__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ net1200 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
X_15888_ clknet_leaf_23_wb_clk_i _02028_ _00696_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14839_ net1207 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
X_08360_ _04034_ _04041_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_3_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16509_ clknet_leaf_1_wb_clk_i _02643_ _01316_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_190_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08291_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__inv_2
XANTENNA__12608__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11323__A2_N net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10212__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12343__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09366__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _06815_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_1
XANTENNA__09905__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
Xfanout325 net328 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_2
Xfanout336 _06994_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
X_09814_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\] net835 net819 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\]
+ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__a221o_1
Xfanout347 _07187_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_2
Xfanout358 net361 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_2
Xfanout369 net373 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1100_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] net695 net840 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout560_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13465__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10279__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\] net830 net826 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\]
+ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08627_ net99 team_02_WB.START_ADDR_VAL_REG\[5\] net955 vssd1 vssd1 vccd1 vccd1 _02633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A _04512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08558_ _03292_ _04226_ _04180_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12518__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ team_02_WB.instance_to_wrap.top.a1.state\[1\] _04184_ net849 net2025 vssd1
+ vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10520_ _04461_ _05963_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nor2_4
XFILLER_0_9_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10451_ _04713_ _04733_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10203__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13170_ _07487_ _07488_ _07501_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nand3b_1
X_10382_ net972 net644 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ net276 net2308 net466 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12253__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10562__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net271 net1901 net472 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__mux2_1
Xhold390 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _06349_ _06512_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_73_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout870 net873 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09109__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15811_ clknet_leaf_10_wb_clk_i _01951_ _00619_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout881 _04538_ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
X_16791_ net1335 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_4
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08686__B team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15742_ clknet_leaf_5_wb_clk_i _01882_ _00550_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12954_ team_02_WB.instance_to_wrap.top.pc\[13\] _06205_ vssd1 vssd1 vccd1 vccd1
+ _07474_ sky130_fd_sc_hd__or2_1
Xhold1090 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11905_ net346 net2551 net486 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
X_15673_ clknet_leaf_124_wb_clk_i _01813_ _00481_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12885_ net506 _05582_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ net1103 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11836_ net352 net1946 net588 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14555_ net1085 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12428__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net354 net2559 net598 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13506_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10718_ _06148_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__and2b_1
X_14486_ net1084 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XANTENNA__10456__B _05061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ net953 _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16225_ clknet_leaf_101_wb_clk_i _02365_ _01033_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13437_ _03036_ _03038_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__xor2_1
X_10649_ _04350_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09596__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11839__Y _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16156_ clknet_leaf_19_wb_clk_i _02296_ _00964_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13368_ net2634 net1018 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[30\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09060__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net1102 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
XANTENNA__12163__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12319_ net282 net2334 net565 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__mux2_1
X_16087_ clknet_leaf_114_wb_clk_i _02227_ _00895_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13299_ team_02_WB.instance_to_wrap.top.pc\[10\] net1054 _06950_ net933 vssd1 vssd1
+ vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13144__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ net1259 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07860_ _03572_ _03582_ _03540_ net329 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_208_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire626_A _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07791_ _03490_ net366 vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__nand2_1
XANTENNA__08596__B net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\] net707 _05045_ _05046_
+ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09520__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09461_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\] net914 net800 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\]
+ _04977_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a221o_1
XFILLER_0_204_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08412_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04106_ vssd1 vssd1 vccd1
+ vccd1 _04120_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09392_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_195_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08343_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12338__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B1 _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout239_A _06424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _03962_ _03988_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13958__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A _05900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12862__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__A_N net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11478__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_2
XANTENNA_fanout775_A _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12801__S _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ _03706_ _03711_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__S net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\] net833 net899 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a22o_1
XANTENNA__09511__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\] net687 net841 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ net353 net1958 net434 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XANTENNA__09411__A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__C _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ net397 _07035_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_120_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12248__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14340_ net1092 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XANTENNA__08672__D team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _05916_ _06110_ _07042_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire512 _05488_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
Xwire523 _05186_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09290__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10503_ _05208_ _05979_ _05978_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_42_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11483_ net411 _06579_ net418 vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14271_ net1108 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16010_ clknet_leaf_37_wb_clk_i _02150_ _00818_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09578__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10434_ net534 _04822_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nor2_1
XANTENNA_input71_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ net623 net938 net1019 net1619 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10563__Y _06080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10365_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] net898 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ _07505_ _07506_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__or2_1
XANTENNA__13126__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12104_ net2306 net358 net582 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_X clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13084_ _06683_ net234 _02860_ net978 _02858_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__o221a_1
X_10296_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] net749 net733 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a221o_1
XANTENNA__11675__X _07161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12035_ net340 net1966 net474 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16774_ net1318 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_13986_ net1124 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
XANTENNA__09502__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15725_ clknet_leaf_49_wb_clk_i _01865_ _00533_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12937_ team_02_WB.instance_to_wrap.top.pc\[23\] _06177_ vssd1 vssd1 vccd1 vccd1
+ _07457_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15656_ clknet_leaf_11_wb_clk_i _01796_ _00464_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12868_ _05742_ _05782_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_199_Right_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14607_ net1222 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_177_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ net284 net2037 net588 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12158__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ clknet_leaf_9_wb_clk_i _01727_ _00395_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ net848 _04355_ _06161_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__nor3_1
XFILLER_0_173_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14538_ net1179 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09281__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14469_ net1172 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XANTENNA__09569__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16208_ clknet_leaf_22_wb_clk_i _02348_ _01016_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16139_ clknet_leaf_16_wb_clk_i _02279_ _00947_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13117__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08792__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08792__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\] net763 net730 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ _03632_ _03633_ _03621_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12621__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ net3 net1033 net989 net1469 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _03561_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3b_1
XFILLER_0_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07774_ net366 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09513_ _05023_ _05025_ _05027_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_88_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13319__A2_N _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12857__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\] net769 _04957_ _04958_
+ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09375_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] net823 net909 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\]
+ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a221o_1
XANTENNA__12068__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08326_ _04015_ _04017_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__nor2_1
XANTENNA__09272__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ _03925_ _03953_ _03960_ _03927_ _03913_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a32o_1
XFILLER_0_201_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08480__B1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08188_ _03888_ _03893_ _03862_ _03868_ _03877_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10383__Y _05900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13200__B _02953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09980__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _05660_ _05662_ _05664_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor4_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\] net832 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\]
+ _05585_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a221o_1
XANTENNA__10840__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ net1147 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XANTENNA__10893__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13771_ net1945 _03265_ net960 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10986__S net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08838__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10839__X _06355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ net999 _06494_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13292__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15510_ clknet_leaf_22_wb_clk_i _01650_ _00318_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15143__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ _06469_ _06500_ _07245_ _06426_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__or4b_1
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ clknet_leaf_66_wb_clk_i net1428 _01298_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XANTENNA__16348__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__C team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15441_ clknet_leaf_2_wb_clk_i _01581_ _00249_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12653_ net285 net2285 net434 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14982__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09799__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11604_ net377 _06940_ _07090_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15372_ clknet_leaf_68_wb_clk_i _01512_ _00185_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_12584_ net277 net2071 net438 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ net1074 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11535_ team_02_WB.instance_to_wrap.top.pc\[6\] _06255_ vssd1 vssd1 vccd1 vccd1 _07027_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07596__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14254_ net1083 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XANTENNA_input74_X net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11466_ _06869_ _06960_ net396 vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13205_ _04732_ net938 net1019 net1514 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a2bb2o_1
X_10417_ _05931_ _05933_ _05335_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__o21a_1
X_14185_ net1231 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
X_11397_ _05931_ _06894_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08979__X _04496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10030__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _07377_ _07414_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__xnor2_1
X_10348_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\] net717 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10279_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\] net926 net796 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\]
+ _05789_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a221o_1
X_13067_ team_02_WB.instance_to_wrap.top.pc\[24\] _07349_ _02845_ _02846_ vssd1 vssd1
+ vccd1 vccd1 _01505_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_146_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ net270 net1932 net477 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16757_ net1301 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XANTENNA__13283__B1 _06759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ net1252 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
XANTENNA__10097__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15708_ clknet_leaf_19_wb_clk_i _01848_ _00516_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ clknet_leaf_71_wb_clk_i _02805_ _01412_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09051__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ clknet_leaf_115_wb_clk_i _01779_ _00447_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10197__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09160_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] net912 net888 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09254__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ _03792_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11597__B1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ net970 net635 net543 vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12616__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08042_ _03721_ _03760_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold901 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10021__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 team_02_WB.instance_to_wrap.top.a1.row1\[15\] vssd1 vssd1 vccd1 vccd1 net2318
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09962__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _05505_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or2_2
Xhold989 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12351__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ _04309_ _04459_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_95_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08875_ net21 net1031 _04432_ net1630 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__o22a_1
X_07826_ _03509_ _03538_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07757_ _03452_ _03477_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout640_A _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A _04379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ _03393_ _03394_ _03377_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09493__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09427_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\] net803 _04930_ _04943_
+ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1170_X net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09358_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\] net772 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a22o_1
XANTENNA__09245__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08309_ _03992_ _04000_ _04007_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10835__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12526__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09289_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\] net924 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ net376 _06606_ _06820_ net383 vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10260__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ _05126_ net657 vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08024__B team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\] net736 net684 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09953__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ _05016_ net387 _06338_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__a21o_1
XANTENNA__11760__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] net767 net751 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__a22o_1
XANTENNA__12261__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ clknet_leaf_21_wb_clk_i _02130_ _00798_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09705__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ net1207 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
X_10064_ _05441_ _05580_ net550 vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__mux2_1
XANTENNA_input34_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__B _06883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_202_Right_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14872_ net1184 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ clknet_leaf_93_wb_clk_i _02730_ _01404_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_13823_ net1138 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08694__B _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10079__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11276__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ clknet_leaf_82_wb_clk_i _00014_ _01349_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13754_ net1832 _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__o21a_1
X_10966_ _06399_ _06478_ net371 vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09484__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10729__B _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ net1004 net1070 _04249_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16473_ clknet_leaf_69_wb_clk_i net1499 _01281_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11291__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13685_ _03200_ _03204_ _03213_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a21oi_1
X_10897_ net667 _06398_ _06407_ net795 _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o221a_1
XFILLER_0_183_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08981__Y _04498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15424_ clknet_leaf_17_wb_clk_i _01564_ _00232_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12636_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] net362 net552 vssd1
+ vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__mux2_1
XANTENNA__09236__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15355_ clknet_leaf_75_wb_clk_i _01495_ _00168_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12436__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ net343 net2336 net443 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11340__S net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ net1129 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XANTENNA__10251__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11518_ team_02_WB.instance_to_wrap.top.pc\[7\] net975 _04347_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__a22o_1
X_15286_ clknet_leaf_84_wb_clk_i _01430_ _00099_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12498_ net337 net2181 net559 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__mux2_1
Xhold208 _02594_ vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold219 team_02_WB.instance_to_wrap.top.a1.row1\[2\] vssd1 vssd1 vccd1 vccd1 net1581
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ net1203 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
X_11449_ _05469_ net663 _06943_ net794 _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o221a_1
XANTENNA__09944__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ net1195 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13119_ _07418_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12171__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14099_ net1072 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XANTENNA__15268__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14887__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ net1061 net1544 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1
+ vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a21o_2
XFILLER_0_163_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ _03331_ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13256__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08591_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09052__Y _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09475__A2 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09212_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] net912 net852 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09227__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09143_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\] net764 net728 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12346__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11103__X _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10242__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] net895 net942 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08025_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] _03746_ _03747_ vssd1 vssd1
+ vccd1 vccd1 _03748_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold720 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1130_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold731 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold742 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09935__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold753 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold797 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10390__A _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12081__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\] net863 net854 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a22o_1
X_08927_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] net958 vssd1 vssd1 vccd1
+ vccd1 _04447_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout855_A _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net167 net1043 net1035 net1383 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_179_Left_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08795__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08910__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07809_ _03512_ _03524_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__a21o_2
XANTENNA__08910__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08789_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04275_ _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10820_ _05061_ _05901_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__C _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09466__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10751_ team_02_WB.instance_to_wrap.top.pc\[25\] team_02_WB.instance_to_wrap.top.pc\[24\]
+ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__and3_1
XFILLER_0_177_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ team_02_WB.START_ADDR_VAL_REG\[10\] net1069 net1002 vssd1 vssd1 vccd1 vccd1
+ net193 sky130_fd_sc_hd__a21o_1
XFILLER_0_48_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10682_ net994 _04419_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12421_ net274 net2000 net457 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__mux2_1
XANTENNA__12256__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14037__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ net1144 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10233__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ net282 net1908 net561 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ _05941_ _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15071_ net1168 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XANTENNA__12780__A _06965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net267 net2174 net571 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XANTENNA__09926__A0 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14022_ net1212 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
X_11234_ net973 _06733_ _06738_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_3_1_0_wb_clk_i_X clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__A0 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ _06669_ _06670_ _06671_ net666 vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\] net889 net869 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__a22o_1
X_11096_ _06542_ _06604_ net371 vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__mux2_1
X_15973_ clknet_leaf_29_wb_clk_i _02113_ _00781_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13486__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14924_ net1215 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
X_10047_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\] net732 _05562_ _05563_
+ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a211o_1
XANTENNA__14500__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 team_02_WB.START_ADDR_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 team_02_WB.instance_to_wrap.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 net1453
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14855_ net1174 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
X_13806_ net1163 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14786_ net1194 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XANTENNA__09457__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ net325 net1869 net481 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16525_ clknet_leaf_0_wb_clk_i _02659_ _01332_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13737_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ _03242_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_158_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10949_ _06141_ _06145_ _06237_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ clknet_leaf_45_wb_clk_i net1450 _01264_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13668_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_80_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09209__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15407_ clknet_leaf_42_wb_clk_i _01547_ _00215_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12619_ net2143 net273 net553 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__mux2_1
XANTENNA__11016__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12166__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16387_ clknet_leaf_89_wb_clk_i _02522_ _01195_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13599_ team_02_WB.instance_to_wrap.top.a1.row1\[58\] _03117_ _03125_ team_02_WB.instance_to_wrap.top.a1.row2\[34\]
+ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10224__A0 _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13275__A1_N _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15338_ clknet_leaf_44_wb_clk_i _01481_ _00151_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15269_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[28\]
+ _00082_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_187_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\] net840 _05342_ _05343_
+ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09047__Y _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\] net818 net884 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_206_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13213__A1_N net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ _04289_ _04311_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__or2_1
X_09692_ net522 _05206_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__and2_1
XANTENNA__09696__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ _03298_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _04272_ sky130_fd_sc_hd__nand2_1
XANTENNA__13229__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_A _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08574_ team_02_WB.instance_to_wrap.top.a1.row1\[58\] _04238_ _04225_ vssd1 vssd1
+ vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09448__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__A1_N net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12865__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13313__X _03006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11007__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout603_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] net926 net812 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a22o_1
XANTENNA__09081__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11963__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\] net782 net746 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09908__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ _03692_ _03703_ _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold550 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] vssd1 vssd1
+ vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold594 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] net778 net682 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ team_02_WB.instance_to_wrap.top.pc\[4\] _05742_ vssd1 vssd1 vccd1 vccd1 _07490_
+ sky130_fd_sc_hd__nand2_1
Xhold1250 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09687__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1261 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ net287 net1775 net482 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1272 team_02_WB.instance_to_wrap.ramload\[30\] vssd1 vssd1 vccd1 vccd1 net2634
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14640_ net1236 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11852_ net274 net2178 net493 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09439__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10803_ net391 _06315_ _06316_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ net1152 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
X_11783_ net288 net1752 net592 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08972__B _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16310_ clknet_leaf_50_wb_clk_i _02450_ _01118_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13522_ _03078_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nor2_1
X_10734_ _04344_ _04349_ _04354_ _04325_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_171_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ clknet_leaf_128_wb_clk_i _02381_ _01049_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13453_ _03038_ _03055_ _02768_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_62_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10665_ team_02_WB.instance_to_wrap.top.pc\[21\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _06182_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10206__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12404_ net355 net1746 net460 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__mux2_1
X_16172_ clknet_leaf_2_wb_clk_i _02312_ _00980_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13384_ team_02_WB.instance_to_wrap.ramload\[13\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[13\] sky130_fd_sc_hd__and2_1
XANTENNA__13089__A2_N net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10596_ _04460_ _04468_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__nand2_4
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09611__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15123_ net1165 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
X_12335_ net339 net2432 net564 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
XANTENNA__15926__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ net1166 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
X_12266_ net325 net2224 net572 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__mux2_1
X_14005_ net1224 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
X_11217_ net374 _06472_ _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__o21a_1
X_12197_ net314 net2480 net578 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11182__A1 _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11148_ net973 _06651_ _06654_ _06655_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15956_ clknet_leaf_3_wb_clk_i _02096_ _00764_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11079_ net953 _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__nand2_1
XANTENNA__09678__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ net1077 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
X_15887_ clknet_leaf_43_wb_clk_i _02027_ _00695_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_201_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14838_ net1083 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14769_ net1229 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16508_ clknet_leaf_6_wb_clk_i _02642_ _01315_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15456__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ _04003_ _04004_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__and2_1
XANTENNA__10996__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16439_ clknet_leaf_42_wb_clk_i net1393 _01247_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_200_Left_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09602__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08810__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12624__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout304 net307 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
Xfanout315 _06914_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
Xfanout326 net328 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_2
Xfanout337 _06994_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_1
X_09813_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\] net921 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a22o_1
XANTENNA__13152__A1_N net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout348 _07187_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
Xfanout359 net361 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_2
X_09744_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\] net735 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\]
+ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a221o_1
XANTENNA__14140__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\] net877 net856 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a22o_1
XANTENNA__08877__B1 _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08626_ net100 net1616 net957 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08629__A0 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08557_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04174_ vssd1 vssd1 vccd1
+ vccd1 _04226_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_120_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08488_ team_02_WB.instance_to_wrap.top.a1.row1\[13\] _04185_ vssd1 vssd1 vccd1 vccd1
+ _02697_ sky130_fd_sc_hd__or2_1
XANTENNA__09841__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15949__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ _04630_ _04652_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__nand2_1
XANTENNA__09054__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] net757 net717 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07604__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _05882_ _05892_ _05895_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__nor4_1
XANTENNA__12534__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14315__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12120_ net283 net1572 net467 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ net263 net2457 net472 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold380 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 team_02_WB.START_ADDR_VAL_REG\[24\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ net414 _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_205_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout860 _04544_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_8
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
X_15810_ clknet_leaf_119_wb_clk_i _01950_ _00618_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_16790_ net1334 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
Xfanout882 _04537_ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_8
Xfanout893 _04533_ vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15741_ clknet_leaf_14_wb_clk_i _01881_ _00549_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12953_ team_02_WB.instance_to_wrap.top.pc\[13\] _06205_ vssd1 vssd1 vccd1 vccd1
+ _07473_ sky130_fd_sc_hd__nand2_1
Xhold1080 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14985__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1091 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net350 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] net486 vssd1
+ vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15672_ clknet_leaf_121_wb_clk_i _01812_ _00480_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12884_ net428 _05627_ _07403_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08983__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14623_ net1126 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XANTENNA__11219__A2 _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11835_ net362 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\] net588 vssd1
+ vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07599__A team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14554_ net1089 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ net358 net1986 net599 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__mux2_1
XANTENNA__09293__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09832__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _06151_ _06233_ _06152_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__o21bai_1
X_14485_ net1257 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _07180_ _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__nor2_2
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16224_ clknet_leaf_18_wb_clk_i _02364_ _01032_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13436_ _03032_ _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__and2_1
XANTENNA__08922__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ _06154_ _06163_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__a21o_1
XANTENNA__09045__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ clknet_leaf_32_wb_clk_i _02295_ _00963_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12444__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ net2510 net1018 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[29\]
+ sky130_fd_sc_hd__and2_1
X_10579_ _04970_ net388 _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__a21o_1
X_15106_ net1079 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12318_ net269 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\] net567 vssd1
+ vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__mux2_1
X_16086_ clknet_leaf_49_wb_clk_i _02226_ _00894_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_184_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13298_ net1632 net982 net964 _02998_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ net1259 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12249_ net257 net2469 net572 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11155__A1 _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap616_A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09899__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15056__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09325__Y _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ _03494_ _03485_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire619_A _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08859__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15939_ clknet_leaf_9_wb_clk_i _02079_ _00747_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11458__A2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09520__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\] net886 net874 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08411_ _04105_ _04111_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__xor2_2
X_09391_ _04886_ _04905_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__nor2_1
XANTENNA__12619__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08342_ _04035_ _04053_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10969__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09823__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ _03962_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09036__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12862__B _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12354__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__B1 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10382__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1210_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13540__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ _03707_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] net817 net907 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\]
+ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a221o_1
XANTENNA__11449__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09658_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] net716 net695 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\]
+ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10121__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ net87 net1566 net955 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_106_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12529__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] net911 net883 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11620_ net1928 net365 net637 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09275__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09814__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _05915_ _06116_ net660 _05691_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_64_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_2
X_10502_ _04950_ _05982_ _05981_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_42_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14270_ net1127 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
Xwire535 _04801_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_2
X_11482_ _05559_ _06006_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ net625 net938 net1019 net1496 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a2bb2o_1
X_10433_ _04865_ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12264__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12582__A0 _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input64_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13152_ net1026 _02917_ net1024 team_02_WB.instance_to_wrap.top.pc\[10\] vssd1 vssd1
+ vccd1 vccd1 _01491_ sky130_fd_sc_hd__a2bb2o_1
X_10364_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] net824 net820 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16277__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12103_ net1685 net344 net582 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
X_13083_ _07427_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__xnor2_1
X_10295_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] net773 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a22o_1
XANTENNA__11137__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12034_ net333 net1800 net475 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__mux2_1
XANTENNA__11688__A2 _07161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 _04397_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_4
X_16773_ net1317 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_13985_ net1258 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ clknet_leaf_2_wb_clk_i _01864_ _00532_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12936_ team_02_WB.instance_to_wrap.top.pc\[24\] _04494_ vssd1 vssd1 vccd1 vccd1
+ _07456_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_124_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08917__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15655_ clknet_leaf_38_wb_clk_i _01795_ _00463_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12439__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ net505 _05671_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11818_ net272 net1871 net589 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
X_14606_ net1075 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
XFILLER_0_201_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08449__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15586_ clknet_leaf_117_wb_clk_i _01726_ _00394_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12798_ _07321_ _07258_ _07247_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__or3b_4
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09805__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14537_ net1221 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11749_ net277 net2389 net596 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13411__X _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ net1092 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16207_ clknet_leaf_43_wb_clk_i _02347_ _01015_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13419_ _03030_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__inv_2
XANTENNA__12174__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14399_ net1115 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XANTENNA__10179__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16138_ clknet_leaf_37_wb_clk_i _02278_ _00946_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09049__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08792__A2 _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13117__A2 _07332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16069_ clknet_leaf_29_wb_clk_i _02209_ _00877_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_08960_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] net771 net758 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a221o_1
X_07911_ _03614_ _03615_ _03617_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08891_ net4 net1029 net986 net1996 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__o22a_1
XFILLER_0_208_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07842_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nand2_1
XANTENNA__10351__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12628__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ _03482_ _03494_ _03495_ _03485_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_142_Left_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09512_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\] net809 net897 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\]
+ _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10103__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\] net713 net838 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\]
+ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a221o_1
XANTENNA__12349__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_A _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09374_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\] net904 net871 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13053__B2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08325_ _04038_ _03321_ net1007 net1668 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_191_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07967__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08256_ _03966_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08480__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _03875_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout885_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] net926 _05584_ _05596_
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_X clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10342__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13770_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\]
+ _03263_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__and3_1
XANTENNA__09496__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _06143_ net652 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] net496
+ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__a221o_1
XANTENNA__13292__B2 _02995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ _06533_ _06566_ _06596_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_179_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12259__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15440_ clknet_leaf_21_wb_clk_i _01580_ _00248_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12652_ net274 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\] net437 vssd1
+ vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__mux2_1
XANTENNA__08683__D team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09248__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ net397 _07016_ net384 vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__o21ai_1
X_15371_ clknet_leaf_68_wb_clk_i _01511_ _00184_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[30\]
+ sky130_fd_sc_hd__dfrtp_2
X_12583_ net283 net2353 net440 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ net1177 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
X_11534_ net670 _07014_ _07025_ net672 _07024_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14253_ net1126 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
X_11465_ _06919_ _06959_ net369 vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13204_ _04691_ net937 net1021 net1443 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10416_ _05378_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14184_ net1111 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
X_11396_ _05381_ _05930_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nor2_1
XANTENNA__09420__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13135_ _07511_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__xnor2_1
X_10347_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] net693 net838 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\]
+ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ _06590_ net234 net231 _02843_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__a2bb2o_1
X_10278_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] _04529_ _05791_ _05792_
+ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__a2111o_1
X_12017_ net262 net2431 net477 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
XANTENNA__08995__X _04512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10333__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16756_ net1300 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_177_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09487__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13283__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ net1252 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15707_ clknet_leaf_29_wb_clk_i _01847_ _00515_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12169__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ _04672_ _06139_ _07355_ _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10478__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16687_ clknet_leaf_70_wb_clk_i _02804_ _01411_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13899_ net1246 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09051__B _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09239__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15638_ clknet_leaf_21_wb_clk_i _01778_ _00446_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10197__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15569_ clknet_leaf_0_wb_clk_i _01709_ _00377_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__X _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _03795_ _03800_ _03815_ _03816_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a22oi_4
XANTENNA__11801__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11597__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09090_ _04593_ _04601_ _04604_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__nor4_1
XFILLER_0_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08041_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03760_ _03761_ vssd1 vssd1
+ vccd1 vccd1 _03763_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_211_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold902 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_2
Xhold924 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12632__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ _05494_ _05496_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__or3_1
Xhold979 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ _04309_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nor2_1
XANTENNA__13496__A_N net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16401__Q team_02_WB.instance_to_wrap.ramload\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout299_A _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ net22 net1030 net987 team_02_WB.instance_to_wrap.ramload\[28\] vssd1 vssd1
+ vccd1 vccd1 _02556_ sky130_fd_sc_hd__o22a_1
XANTENNA__10324__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1006_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _03536_ _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__and2_1
XANTENNA__09190__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12868__A _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07756_ _03449_ _03451_ _03477_ _03445_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__a31o_1
XFILLER_0_189_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07687_ _03403_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__nand2_1
XANTENNA__12079__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\] net834 net920 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\]
+ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09357_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] net783 net719 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12807__S _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11711__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12785__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _04020_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09288_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] net887 net867 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08239_ _03942_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11250_ net421 _06749_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nand2_1
XANTENNA__09402__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10201_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\] net752 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__a22o_1
XANTENNA__08024__C team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11181_ _05041_ _05945_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12542__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14323__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _05647_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13501__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14940_ net1199 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
X_10063_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] _04330_ net648 team_02_WB.instance_to_wrap.top.a1.instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a22o_1
XANTENNA__09181__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ net1186 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
X_16610_ clknet_leaf_96_wb_clk_i _02729_ _01403_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13822_ net1147 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
XANTENNA__09469__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13753_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] _03254_ net950 vssd1
+ vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ clknet_leaf_84_wb_clk_i _00013_ _01348_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10965_ _06076_ _06079_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14993__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ net348 net2077 net430 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13684_ net1381 _03199_ net1066 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__o21ai_1
X_16472_ clknet_leaf_71_wb_clk_i net1520 _01280_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
X_10896_ net656 _06402_ _06409_ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__o211a_1
X_15423_ clknet_leaf_62_wb_clk_i _01563_ _00231_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ net1666 net355 net554 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__mux2_1
XANTENNA__10585__X _06102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11579__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15354_ clknet_leaf_76_wb_clk_i _01494_ _00167_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12566_ net338 net1997 net442 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09641__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14305_ net1256 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11517_ net1000 _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nor2_1
X_15285_ clknet_leaf_70_wb_clk_i _01429_ _00098_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ net326 net1818 net557 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold209 team_02_WB.instance_to_wrap.ramstore\[16\] vssd1 vssd1 vccd1 vccd1 net1571
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ net1199 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
X_11448_ _05465_ net660 _06116_ _05466_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12960__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14167_ net1185 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XANTENNA__12452__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ net421 _06037_ _06388_ _06110_ _06014_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a32o_1
XANTENNA__08869__C net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ _07372_ _07373_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__and2b_1
X_14098_ net1177 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13049_ net1027 _02831_ net1024 team_02_WB.instance_to_wrap.top.pc\[27\] vssd1 vssd1
+ vccd1 vccd1 _01508_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_56_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10306__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__buf_4
XANTENNA__09172__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07610_ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] _03324_ _03328_ vssd1 vssd1
+ vccd1 vccd1 _03333_ sky130_fd_sc_hd__and3_1
X_08590_ net70 net69 net41 net40 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_85_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16739_ net1284 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_163_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09997__A _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] net867 _04715_ _04727_
+ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12627__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\] net736 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09632__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] net819 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08024_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] team_02_WB.instance_to_wrap.top.a1.dataIn\[6\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold710 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold743 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12362__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15212__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] net894 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a22o_1
XANTENNA__10390__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout583_A _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ net1421 _04446_ net930 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XANTENNA__09699__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09163__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ net168 net1042 net1034 net1470 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout750_A _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ _03530_ _03527_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2b_1
X_08788_ net1060 net648 _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a21o_2
XANTENNA__12748__D _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _03422_ _03459_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10750_ team_02_WB.instance_to_wrap.top.pc\[23\] _06266_ vssd1 vssd1 vccd1 vccd1
+ _06267_ sky130_fd_sc_hd__and2_1
XANTENNA__09871__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09409_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\] net763 _04923_ _04924_
+ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_164_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ team_02_WB.instance_to_wrap.top.pc\[14\] _06197_ vssd1 vssd1 vccd1 vccd1
+ _06198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ net289 net1783 net455 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ net269 net2256 net562 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15210__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _05212_ _05940_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__nor2_1
X_15070_ net1247 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
X_12282_ net258 net2221 net568 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14021_ net1176 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
X_11233_ _06186_ net653 _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10581__A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ net379 _06396_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] _04529_ net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a22o_1
X_15972_ clknet_leaf_36_wb_clk_i _02112_ _00780_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11095_ _06072_ _06098_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__or2_1
XANTENNA__08986__A team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14923_ net1124 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
X_10046_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\] net705 net685 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_203_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold70 _02623_ vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_02_WB.instance_to_wrap.ramstore\[28\] vssd1 vssd1 vccd1 vccd1 net1443
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 _02585_ vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ net1205 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13805_ net1164 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__inv_2
X_14785_ net1260 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
X_11997_ net321 net2590 net478 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16524_ clknet_leaf_127_wb_clk_i _02658_ _01331_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13736_ _03244_ net951 _03243_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__and3b_1
X_10948_ _06140_ net652 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] net497
+ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16455_ clknet_leaf_44_wb_clk_i net1444 _01263_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10879_ _06066_ _06090_ net369 vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__mux2_1
XANTENNA__12447__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_80_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15406_ clknet_leaf_45_wb_clk_i _01546_ _00214_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12618_ net1682 net291 net552 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ team_02_WB.instance_to_wrap.top.a1.row1\[114\] _03121_ _03123_ team_02_WB.instance_to_wrap.top.a1.row2\[42\]
+ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__a22o_1
X_16386_ clknet_leaf_89_wb_clk_i _02521_ _01194_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09614__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10224__A1 _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08968__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15337_ clknet_leaf_44_wb_clk_i _01480_ _00150_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12549_ net271 net1529 net445 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_max_cap646_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15235__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_1 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[27\]
+ _00081_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_14219_ net1137 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XANTENNA__12182__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15199_ net1245 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09393__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\] net920 net810 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_206_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ team_02_WB.instance_to_wrap.top.a1.instruction\[5\] _04309_ _04339_ _04316_
+ _04268_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__o32a_1
XANTENNA__09145__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _05187_ _05206_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__and2_1
Xfanout1090 net1094 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
X_08642_ net1059 _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13229__B2 _05760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10160__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ team_02_WB.instance_to_wrap.top.a1.halfData\[0\] _04228_ _04230_ _02812_
+ _04227_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12865__B _05491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A _07013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12357__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1073_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09605__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09125_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\] _04641_ vssd1 vssd1 vccd1
+ vccd1 _04642_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08959__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09056_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\] net763 _04570_ _04572_
+ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout798_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _03703_ _03691_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__and2b_1
XANTENNA__12092__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09238__Y _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold551 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold562 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold584 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\] net734 net839 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a22o_1
X_08909_ net1445 _04436_ net930 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XANTENNA__11479__B1 _06833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\] net804 net882 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ _05401_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1
+ net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ net274 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\] net485 vssd1
+ vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
Xhold1262 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1273 team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net2635
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11851_ net290 net2089 net491 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ net391 _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nor2_1
X_14570_ net1176 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
X_11782_ net278 net2053 net592 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09844__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10733_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _06161_ _06248_ net953 vssd1
+ vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a31o_1
X_13521_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[1\] team_02_WB.instance_to_wrap.top.pad.keyCode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__or4b_2
XANTENNA__12267__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13452_ _02764_ _02765_ _03036_ _02763_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__or4_1
X_16240_ clknet_leaf_26_wb_clk_i _02380_ _01048_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input94_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10664_ team_02_WB.instance_to_wrap.top.pc\[21\] _06180_ vssd1 vssd1 vccd1 vccd1
+ _06181_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12403_ net359 net2145 net461 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__mux2_1
X_13383_ team_02_WB.instance_to_wrap.ramload\[12\] net1013 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[12\] sky130_fd_sc_hd__and2_1
X_16171_ clknet_leaf_15_wb_clk_i _02311_ _00979_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12791__A _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10595_ _04460_ _04468_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_153_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09429__X _04946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12334_ net332 net2350 net564 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__mux2_1
X_15122_ net1165 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15053_ net1164 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
X_12265_ net321 net1830 net572 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11613__A2_N net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ net1238 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
X_11216_ net422 _06475_ _06638_ _06471_ net377 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__a221o_1
XANTENNA__09375__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net306 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] net579 vssd1
+ vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11147_ _06177_ net653 net494 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] net496
+ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09127__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11078_ _06580_ _06584_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__a21oi_4
X_15955_ clknet_leaf_56_wb_clk_i _02095_ _00763_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10029_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\] net815 net798 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__a221o_1
X_14906_ net1089 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
X_15886_ clknet_leaf_46_wb_clk_i _02026_ _00694_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08886__B2 net2477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14837_ net1242 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_201_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14768_ net1226 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09835__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16507_ clknet_leaf_6_wb_clk_i _02641_ _01314_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13719_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__or2_1
X_14699_ net1120 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16183__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16438_ clknet_leaf_83_wb_clk_i net1497 _01246_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16369_ clknet_leaf_128_wb_clk_i _02509_ _01177_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09366__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 net307 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08574__A0 team_02_WB.instance_to_wrap.top.a1.row1\[58\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09812_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] net823 net853 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\]
+ _05316_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__a221o_1
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
XANTENNA__12640__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
Xfanout349 _07187_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_1
XFILLER_0_185_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09118__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] net779 net775 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout281_A _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout379_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\] net913 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\]
+ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_19_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08877__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10133__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ net101 net1589 net956 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1190_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__A _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _04489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08556_ net1047 _04183_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_120_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09826__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_147_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12087__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _04168_ _04179_ _04183_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout713_A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1243_X net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\] net749 net721 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a221o_1
XANTENNA__13500__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\] net832 net894 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\]
+ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09039_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] net887 net876 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\]
+ _04553_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09357__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ net267 net2569 net471 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold370 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ net398 _06346_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__o21a_1
Xhold392 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__Y _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 _04544_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
XANTENNA__09109__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
XFILLER_0_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout883 _04537_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 net897 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_8
X_15740_ clknet_leaf_20_wb_clk_i _01880_ _00548_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12952_ team_02_WB.instance_to_wrap.top.pc\[14\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _07472_ sky130_fd_sc_hd__nand2_1
Xhold1070 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ net364 net2135 net486 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
Xhold1092 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15671_ clknet_leaf_115_wb_clk_i _01811_ _00479_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12883_ _07387_ _07401_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_64_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ net1191 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
X_11834_ net354 net1797 net590 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14553_ net1093 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
XANTENNA__07599__B team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11765_ net342 net1988 net597 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_200_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13504_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__or4_1
X_10716_ team_02_WB.instance_to_wrap.top.pc\[24\] _06172_ _06232_ vssd1 vssd1 vccd1
+ vccd1 _06233_ sky130_fd_sc_hd__a21oi_1
XANTENNA_input97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11696_ _04458_ _04468_ _07177_ _07181_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14484_ net1238 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16223_ clknet_leaf_59_wb_clk_i _02363_ _01031_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13435_ _03030_ _02765_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__or2_1
X_10647_ _04344_ _04349_ _06161_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__and3_1
XANTENNA__13212__A1_N net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ team_02_WB.instance_to_wrap.ramload\[28\] net1018 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[28\] sky130_fd_sc_hd__and2_1
X_16154_ clknet_leaf_18_wb_clk_i _02294_ _00962_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10578_ _05017_ net388 vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15105_ net1074 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
X_12317_ net261 net2349 net565 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__mux2_1
X_16085_ clknet_leaf_40_wb_clk_i _02225_ _00893_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13297_ team_02_WB.instance_to_wrap.top.pc\[11\] net1053 _06931_ net935 vssd1 vssd1
+ vccd1 vccd1 _02998_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_197_Left_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08998__X _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15036_ net1228 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
XANTENNA__13227__A1_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ net249 net1694 net574 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13144__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_max_cap511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ net246 net2195 net579 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14241__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15938_ clknet_leaf_118_wb_clk_i _02078_ _00746_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10115__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09520__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15869_ clknet_leaf_12_wb_clk_i _02009_ _00677_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08410_ _04105_ _04111_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nand2b_1
X_09390_ _04886_ _04905_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08341_ _04030_ _04040_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08272_ _03981_ _03986_ _03964_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a21o_2
XFILLER_0_144_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12635__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09587__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1036_A _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09339__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__X _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16079__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07987_ _03645_ _03695_ _03696_ net256 vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout663_A _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09726_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\] net893 net869 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09511__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] net776 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11714__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08608_ net88 net1753 _04261_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
X_09588_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] net820 net870 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _03313_ _04184_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ net384 _06382_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__nand2_1
XANTENNA__11082__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire503 _05735_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10501_ _05985_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__nor2_1
Xwire514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_174_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_2
X_11481_ net1693 net325 net638 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XANTENNA__12545__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_2
Xwire547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_2
X_13220_ _05375_ net936 net1020 net1392 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a2bb2o_1
X_10432_ _04907_ _05948_ _04908_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09578__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13151_ _06952_ net233 _02916_ net977 _02915_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__o221a_1
X_10363_ net368 _05876_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ net1822 net341 net581 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
X_13082_ _04970_ _06180_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__xnor2_1
X_10294_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] net681 net677 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\]
+ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a221o_1
XANTENNA_input57_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ net336 net1802 net477 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__mux2_1
XANTENNA__12280__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout680 _04407_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_4
XANTENNA__15307__D team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout691 _04397_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_16772_ net1316 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
X_13984_ net1103 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_189_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15723_ clknet_leaf_114_wb_clk_i _01863_ _00531_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09502__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12935_ team_02_WB.instance_to_wrap.top.pc\[24\] _04491_ _04493_ vssd1 vssd1 vccd1
+ vccd1 _07455_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15654_ clknet_leaf_7_wb_clk_i _01794_ _00462_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ net506 _05582_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14605_ net1126 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
X_11817_ net291 net2423 net588 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ clknet_leaf_100_wb_clk_i _01725_ _00393_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12797_ _07311_ _07312_ _07320_ _07306_ _07294_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_32_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14536_ net1104 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
X_11748_ net282 net2503 net598 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
XANTENNA__08933__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14467_ net1134 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XANTENNA__12455__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _07163_ _07164_ _06021_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a21o_1
XFILLER_0_181_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16206_ clknet_leaf_45_wb_clk_i _02346_ _01014_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13418_ net1066 _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nand2_1
XANTENNA__09569__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14398_ net1190 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_180_Right_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16137_ clknet_leaf_111_wb_clk_i _02277_ _00945_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09049__B _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ net2636 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[11\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16068_ clknet_leaf_32_wb_clk_i _02208_ _00876_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12190__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _03571_ _03601_ _03626_ _03605_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__or4b_1
X_15019_ net1167 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
X_08890_ net5 net1029 net986 net2410 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__o22a_1
XANTENNA__10336__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire631_A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ _03517_ _03521_ _03523_ _03553_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__or4_1
XANTENNA__09741__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _03448_ _03460_ _03483_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__and3_1
XANTENNA_wire517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\] net825 net919 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09071__Y _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\] net777 net842 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09373_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\] net835 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\]
+ _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08324_ _04031_ _04036_ _04014_ _04017_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o2bb2a_1
X_08255_ _03947_ _03967_ _03968_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__or3_1
XANTENNA__12365__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1153_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08186_ _03888_ _03893_ _03862_ _03871_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15469__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09980__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout878_A _04538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11709__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1206_X net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09193__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11827__A0 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\] net786 _05224_ _05225_
+ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__a211o_1
X_10981_ team_02_WB.instance_to_wrap.top.pc\[27\] _06269_ vssd1 vssd1 vccd1 vccd1
+ _06494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13292__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _07243_ _06687_ _06658_ _06627_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12651_ net288 net1762 net435 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__mux2_1
XANTENNA__15213__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08066__A1_N _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ net389 _07089_ _07088_ net395 vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__o211a_1
XANTENNA__09799__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _06626_ net2513 net441 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15370_ clknet_leaf_68_wb_clk_i _01510_ _00183_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[29\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08980__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14321_ net1221 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ _05649_ _05917_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12275__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252_ net1214 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
X_11464_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08759__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13203_ net1545 net1021 net939 _04650_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__a22o_1
X_10415_ net519 _05334_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11395_ _06013_ _06892_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__nor2_1
X_14183_ net1181 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16394__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10030__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] net685 net842 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a22o_1
X_13134_ _07476_ _07478_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__nand2_1
XANTENNA__09971__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ net978 _07432_ _02844_ _07337_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__o31ai_1
X_10277_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\] net820 net898 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\]
+ _05793_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__a221o_1
XANTENNA__12858__A2 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09184__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ net268 net2437 net476 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12798__X _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11530__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16755_ net1299 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
X_13967_ net1248 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XANTENNA__13283__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10097__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ clknet_leaf_53_wb_clk_i _01846_ _00514_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12918_ _07356_ _07436_ _07357_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__o21a_1
XANTENNA__08695__C1 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16686_ clknet_leaf_71_wb_clk_i _02803_ _01410_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13898_ net1246 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_192_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15637_ clknet_leaf_31_wb_clk_i _01777_ _00445_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12849_ _06190_ net526 vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_201_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ clknet_leaf_23_wb_clk_i _01708_ _00376_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14519_ net1185 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XANTENNA__12185__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15499_ clknet_leaf_113_wb_clk_i _01639_ _00307_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _03760_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_211_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold903 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold914 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold936 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09962__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold969 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] net883 _05492_ _05507_
+ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a211o_1
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08942_ _04270_ _04288_ _04318_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__and3_2
XANTENNA__09175__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ net23 net1030 net987 net2633 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__o22a_1
XANTENNA__08130__C _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ _03510_ _03534_ _03502_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09523__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07755_ _03449_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout361_A _07069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13274__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout459_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__X _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07686_ _03406_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__nor2_1
XANTENNA__11285__B2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09425_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\] net826 net908 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\] net752 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\]
+ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XFILLER_0_191_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _03997_ _04018_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12095__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09287_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\] _04529_ net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1156_X net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08238_ _03914_ _03927_ _03905_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10260__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08169_ _03865_ _03867_ _03876_ _03882_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__o311a_2
X_10200_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\] net759 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10012__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11180_ net1675 net277 net637 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XANTENNA__09953__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ net428 _05646_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__and2_1
XANTENNA__09166__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ net506 vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__inv_2
XANTENNA__09705__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__A3 _04346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11512__A2 _07001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ net1107 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XANTENNA__12778__B _06902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09433__A _04928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ net1150 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10079__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16540_ clknet_leaf_86_wb_clk_i _02667_ _01347_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[63\]
+ sky130_fd_sc_hd__dfstp_1
X_13752_ _03254_ net950 _03253_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__and3b_1
X_10964_ net377 _06475_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12703_ net352 net1785 net430 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16471_ clknet_leaf_83_wb_clk_i net1608 _01279_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13683_ _03206_ _03212_ net1141 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a21oi_1
X_10895_ _06122_ _06357_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11902__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15422_ clknet_leaf_4_wb_clk_i _01562_ _00230_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12634_ net1886 net358 net553 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15353_ clknet_leaf_78_wb_clk_i _01493_ _00166_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12565_ net330 net2564 net442 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ net1081 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10251__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ _06256_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__or2_1
X_15284_ clknet_leaf_67_wb_clk_i _01428_ _00097_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ net321 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\] net556 vssd1
+ vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ net1085 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
X_11447_ net420 _06514_ _06941_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10003__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09608__A _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ _05932_ net662 net659 _05335_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__a22o_1
XANTENNA__09944__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14166_ net1096 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10329_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__a22o_1
XANTENNA__16502__Q team_02_WB.START_ADDR_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ net790 _07332_ _07515_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__a211o_1
X_14097_ net1229 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
XANTENNA__09157__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ _06494_ net235 _02828_ net977 _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1250 net1252 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_4
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_4
XFILLER_0_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13256__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14999_ net1133 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16738_ net1283 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_76_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16669_ clknet_leaf_66_wb_clk_i _02786_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11812__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\] net826 net806 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\]
+ _04726_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09141_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] net739 net723 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\]
+ _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11414__A1_N net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__inv_2
X_08023_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] team_02_WB.instance_to_wrap.top.a1.dataIn\[2\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] team_02_WB.instance_to_wrap.top.a1.dataIn\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__or4_2
Xhold700 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12643__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold711 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold733 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold744 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold766 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold799 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net791 net650 _05490_
+ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout1116_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] net1009 _04444_ _04445_ vssd1
+ vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a22o_1
XANTENNA__12879__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A _07214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ net1583 net1044 net1036 net1475 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ _03484_ _03528_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08787_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] net997 _04329_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout743_A _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _03443_ _03447_ _03452_ _03457_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a311o_4
XTAP_TAPCELL_ROW_0_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout910_A _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07669_ _03345_ net949 _03361_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_165_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11722__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\] net703 net683 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10481__A2 _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ net789 _05740_ _06127_ _06196_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__o22a_2
XFILLER_0_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\] net798 _04843_ _04855_
+ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11023__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12350_ net261 net2093 net562 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07634__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10233__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ _06584_ _06798_ _06802_ _06037_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12281_ net250 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] net571 vssd1
+ vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XANTENNA__12553__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ net1099 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
X_11232_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] net495 _06736_ net1001 net497
+ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__a221o_1
XANTENNA__13183__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13183__B2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10581__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ net374 _06386_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09139__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\] net923 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a22o_1
X_11094_ _05983_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__xnor2_1
X_15971_ clknet_leaf_27_wb_clk_i _02111_ _00779_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12789__A _06344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13486__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12694__A0 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\] net770 net694 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__a22o_1
X_14922_ net1179 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
Xhold60 team_02_WB.instance_to_wrap.ramstore\[21\] vssd1 vssd1 vccd1 vccd1 net1422
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_02_WB.START_ADDR_VAL_REG\[22\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 _02590_ vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14853_ net1117 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold93 team_02_WB.instance_to_wrap.top.a1.row1\[115\] vssd1 vssd1 vccd1 vccd1 net1455
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ net1366 _03288_ net960 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__o21a_1
X_14784_ net1080 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11996_ net317 net2494 net478 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09311__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08325__A2_N _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16523_ clknet_leaf_6_wb_clk_i _02657_ _01330_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13735_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ _03240_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10947_ net999 _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_158_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16454_ clknet_leaf_71_wb_clk_i net1515 _01262_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13666_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\] _03199_ vssd1 vssd1 vccd1
+ vccd1 _03200_ sky130_fd_sc_hd__and2_1
X_10878_ net396 _06390_ net383 vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15405_ clknet_leaf_48_wb_clk_i _01545_ _00213_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12617_ net2493 net276 net552 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16385_ clknet_leaf_89_wb_clk_i _02520_ _01193_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13597_ team_02_WB.instance_to_wrap.top.a1.row2\[18\] _03124_ _03126_ team_02_WB.instance_to_wrap.top.a1.row2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15336_ clknet_leaf_44_wb_clk_i _01479_ _00149_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12548_ net263 net2465 net445 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12971__B _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12463__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15267_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[26\]
+ _00080_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net250 net2031 net558 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__mux2_1
XANTENNA__09378__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14218_ net1127 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
X_15198_ net1245 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
X_14149_ net1172 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_169_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11807__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _04278_ _04289_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nand2_2
X_09690_ net522 _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1080 net1081 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_4
XANTENNA__09550__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1091 net1093 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_4
X_08641_ team_02_WB.instance_to_wrap.top.a1.instruction\[14\] net1060 vssd1 vssd1
+ vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand2b_1
XANTENNA__13229__A2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ net2522 _04236_ _04225_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XANTENNA__09302__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12638__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10947__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09605__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_A _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1066_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10215__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09124_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] net897 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a22o_1
XANTENNA__09947__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09081__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09055_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] net683 net678 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a22o_1
XANTENNA__12373__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14154__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08006_ _03648_ _03690_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__or2_1
XANTENNA__09908__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold541 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout693_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold552 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold574 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1119_X net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] net774 _05472_ _05473_
+ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_5_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ net1047 _04193_ _04205_ net1009 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a32o_1
XANTENNA__11479__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09888_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\] net828 net824 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a221o_1
Xhold1230 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ net156 net1042 net1034 net1388 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
Xhold1263 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 team_02_WB.instance_to_wrap.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net2636
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ net277 net2321 net490 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
X_10801_ _04589_ net405 vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nor2_1
XANTENNA__12548__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_X net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net282 net2482 net594 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[5\] team_02_WB.instance_to_wrap.top.pad.keyCode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__or4b_2
X_10732_ _04349_ _04354_ _04344_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13451_ _02765_ _03049_ _03054_ _03041_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15221__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10663_ _06128_ _06179_ _04490_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12402_ net342 net2372 net459 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__mux2_1
X_16170_ clknet_leaf_38_wb_clk_i _02310_ _00978_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10206__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ _04462_ _06109_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__or2_2
X_13382_ net2637 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[11\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_input87_A wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15121_ net1162 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
X_12333_ net334 net1955 net565 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12283__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ net1230 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
X_12264_ net317 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\] net572 vssd1
+ vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14003_ net1078 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
X_11215_ net418 _06719_ _06355_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12195_ net299 net2369 net578 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
XANTENNA__09780__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15822__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_X net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ net998 _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11077_ net672 _06566_ _06585_ net671 _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__a221o_2
X_15954_ clknet_leaf_55_wb_clk_i _02094_ _00762_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10028_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\] net827 net921 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__a22o_1
XANTENNA__09532__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ net1098 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
X_15885_ clknet_leaf_40_wb_clk_i _02025_ _00693_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14836_ net1194 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_201_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12966__B _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ net1220 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12458__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ net252 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\] net479 vssd1
+ vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
X_16506_ clknet_leaf_0_wb_clk_i _02640_ _01313_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13718_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\] net950 vssd1 vssd1 vccd1
+ vccd1 _02769_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14698_ net1178 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16437_ clknet_leaf_71_wb_clk_i net1468 _01245_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
X_13649_ net1068 net1010 _07339_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16368_ clknet_leaf_25_wb_clk_i _02508_ _01176_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09063__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15319_ clknet_leaf_83_wb_clk_i _01462_ _00132_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12193__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16299_ clknet_leaf_114_wb_clk_i _02439_ _01107_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10905__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_1
X_09811_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] net861 _05315_ _05327_
+ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__a211o_1
Xfanout317 net320 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09771__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout328 _06975_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
XANTENNA_wire547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout339 net341 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlymetal6s2s_1
X_16785__1329 vssd1 vssd1 vccd1 vccd1 _16785__1329/HI net1329 sky130_fd_sc_hd__conb_1
XFILLER_0_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09742_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\] net683 _05256_ _05257_
+ _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11109__Y _06618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] net928 net861 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08877__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08624_ net102 team_02_WB.START_ADDR_VAL_REG\[8\] net955 vssd1 vssd1 vccd1 vccd1
+ _02636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08555_ _04220_ _04221_ _04224_ net793 net1494 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout441_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12368__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1183_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_194_Right_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08486_ _04168_ _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09054__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\] net745 net685 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1236_X net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__A1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\] net810 net864 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ _04547_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14612__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net398 _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__nand2_1
Xhold393 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _04403_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_8
Xfanout851 _03195_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_2
Xfanout862 _04543_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_8
Xfanout873 _04540_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
Xfanout884 _04537_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09514__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 net897 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_8
X_12951_ team_02_WB.instance_to_wrap.top.pc\[14\] _06200_ vssd1 vssd1 vccd1 vccd1
+ _07471_ sky130_fd_sc_hd__nor2_1
XANTENNA__15216__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1071 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13662__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ net354 net2488 net487 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__mux2_1
Xhold1082 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
X_15670_ clknet_leaf_22_wb_clk_i _01810_ _00478_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1093 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net427 _05627_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__xnor2_1
X_14621_ net1206 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ net360 net2599 net589 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14552_ net1195 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11764_ net339 net1967 net596 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09293__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13503_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16717__1276 vssd1 vssd1 vccd1 vccd1 _16717__1276/HI net1276 sky130_fd_sc_hd__conb_1
XFILLER_0_165_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10715_ _06231_ _06173_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and2b_1
XFILLER_0_193_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14483_ net1080 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
X_11695_ _04569_ _07138_ _07174_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11910__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ clknet_leaf_5_wb_clk_i _02362_ _01030_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13434_ _03036_ _02767_ _02768_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ net848 _06161_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__nand2_1
XANTENNA__10593__Y _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ clknet_leaf_123_wb_clk_i _02293_ _00961_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13365_ net1630 net1018 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[27\]
+ sky130_fd_sc_hd__and2_1
X_10577_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_51_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08504__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ net1072 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XANTENNA__10060__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net265 net2205 net566 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16084_ clknet_leaf_123_wb_clk_i _02224_ _00892_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ net1983 net982 net964 _02997_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__a22o_1
X_15035_ net1230 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
X_12247_ net254 net1739 net573 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12178_ net243 net1993 net578 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16000__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ net418 _06636_ _06355_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__o21a_1
XANTENNA_max_cap504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13301__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15937_ clknet_leaf_100_wb_clk_i _02077_ _00745_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08859__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15868_ clknet_leaf_19_wb_clk_i _02008_ _00676_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16150__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14819_ net1132 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XANTENNA_wire507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12188__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__B1 _07337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799_ clknet_leaf_115_wb_clk_i _01939_ _00607_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11615__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _04040_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08271_ _03981_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09036__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__B1 _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07598__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10051__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12651__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13540__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ _03696_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\] _04529_ _04530_
+ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\] _05241_ vssd1 vssd1 vccd1
+ vccd1 _05242_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09656_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\] net684 _05171_ _05172_
+ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09261__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ net89 net1512 net956 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XANTENNA__12098__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout823_A _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\] net894 net940 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _04222_ net1655 _04186_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09275__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__nor2_1
XANTENNA__11730__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_2
X_11480_ _06837_ _06974_ _06971_ net604 vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_2
X_10431_ _04951_ _05947_ _04948_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_150_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09983__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ _07383_ _07411_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__xnor2_1
X_10362_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12101_ net2006 net330 net580 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XANTENNA__12561__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\] net769 net721 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a22o_1
X_13081_ net231 _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__nand2_1
X_12032_ net325 net1952 net474 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
Xhold190 team_02_WB.instance_to_wrap.ramload\[17\] vssd1 vssd1 vccd1 vccd1 net1552
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _05964_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 _04402_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_4
X_16771_ net1315 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
Xfanout692 _04397_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13983_ net1108 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XANTENNA__13295__B1 _06908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15722_ clknet_leaf_32_wb_clk_i _01862_ _00530_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11905__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ team_02_WB.instance_to_wrap.top.pc\[25\] _06171_ vssd1 vssd1 vccd1 vccd1
+ _07454_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_161_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15653_ clknet_leaf_26_wb_clk_i _01793_ _00461_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ _05489_ _05491_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14604_ net1215 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_1_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11816_ net276 net2297 net588 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ clknet_leaf_110_wb_clk_i _01724_ _00392_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12796_ _07313_ _07315_ _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_194_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535_ net1180 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
X_11747_ net270 net2577 net599 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11640__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16784__1328 vssd1 vssd1 vccd1 vccd1 _16784__1328/HI net1328 sky130_fd_sc_hd__conb_1
XANTENNA__13421__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10281__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ net1130 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
X_11678_ _05016_ _05037_ _05972_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ clknet_leaf_50_wb_clk_i _02345_ _01013_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13417_ team_02_WB.instance_to_wrap.top.lcd.currentState\[1\] net1052 net962 vssd1
+ vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] net995 vssd1 vssd1 vccd1
+ vccd1 _06146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14397_ net1181 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10033__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09974__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ clknet_leaf_11_wb_clk_i _02276_ _00944_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ net1469 net1016 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[10\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_122_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12471__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16067_ clknet_leaf_27_wb_clk_i _02207_ _00875_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap621_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13279_ team_02_WB.instance_to_wrap.top.pc\[20\] team_02_WB.instance_to_wrap.top.ru.state\[5\]
+ _06705_ net935 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a22o_1
XANTENNA__09346__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ net1155 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XANTENNA__09726__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _03521_ _03523_ _03553_ _03517_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__o31ai_1
X_07771_ _03474_ _03489_ _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13286__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15083__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\] net829 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\]
+ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__a221o_1
XANTENNA__16666__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09441_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\] net781 net745 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\] net916 net865 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10020__A _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08323_ _04031_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12646__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11403__X _06901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08254_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10674__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16415__Q team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13210__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ _03901_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout404_A _05900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1146_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10024__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10575__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12381__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716__1275 vssd1 vssd1 vccd1 vccd1 _16716__1275/HI net1275 sky130_fd_sc_hd__conb_1
XANTENNA_fanout1101_X net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07969_ _03690_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout940_A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__B1 _06679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13211__A1_N _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\] net750 net734 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a22o_1
X_10980_ _06236_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_74_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09496__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09639_ _05149_ _05151_ _05153_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__or4_1
XANTENNA__11551__A2_N _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12650_ net278 net2403 net434 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__mux2_1
XANTENNA_input104_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13226__A1_N net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11601_ net498 net385 _06289_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a21boi_1
X_12581_ net264 net2518 net441 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__mux2_1
XANTENNA__12556__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11460__S net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14320_ net1226 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11313__X _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13241__A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11532_ net654 _07019_ _07023_ net794 _07022_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_135_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ net1125 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
X_11463_ _05514_ net657 _06113_ _05512_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_151_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13202_ net635 net936 net1020 net1386 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10414_ _05381_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09956__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14182_ net1212 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XANTENNA__10566__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11394_ _05380_ _06012_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09420__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11696__A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15168__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13133_ net1026 _02901_ net1023 team_02_WB.instance_to_wrap.top.pc\[13\] vssd1 vssd1
+ vccd1 vccd1 _01494_ sky130_fd_sc_hd__a2bb2o_1
X_10345_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\] net733 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12291__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09708__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _07360_ _07431_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nor2_1
X_10276_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] net906 net886 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ net257 net2003 net474 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XANTENNA__14800__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08931__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10599__X _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16754_ net1298 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_13966_ net1248 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
XANTENNA__09487__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15705_ clknet_leaf_125_wb_clk_i _01845_ _00513_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12917_ _07356_ _07436_ _07357_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__o21ai_1
X_16685_ clknet_leaf_65_wb_clk_i _02802_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_13897_ net1244 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15636_ clknet_leaf_3_wb_clk_i _01776_ _00444_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ net531 _06188_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__xor2_1
XANTENNA__09239__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__B _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ clknet_leaf_46_wb_clk_i _01707_ _00375_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12466__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ _07019_ _07095_ _07112_ _07136_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_83_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14518_ net1106 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10254__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15498_ clknet_leaf_38_wb_clk_i _01638_ _00306_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14449_ net1222 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__A0 _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold904 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold915 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold926 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16119_ clknet_leaf_114_wb_clk_i _02259_ _00927_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold937 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_max_cap624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold959 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\] net829 net859 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\]
+ _05506_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08941_ _04336_ _04457_ _04309_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_209_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09175__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ net25 net1032 net988 net2344 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_209_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07823_ _03544_ _03545_ _03540_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07754_ _03461_ _03462_ _03443_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__a21boi_2
XANTENNA__07592__D_N team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ _03363_ _03395_ _03404_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout354_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _04935_ _04937_ _04938_ _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09355_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] net743 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a22o_1
XANTENNA__13431__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12376__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1263_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09286_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\] net876 net860 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ _03823_ _03926_ _03951_ _03911_ _03924_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o2111ai_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09938__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ _03880_ _03883_ _03885_ _03879_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__o22a_1
XANTENNA__09402__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09257__Y _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03762_ _03796_ vssd1 vssd1
+ vccd1 vccd1 _03819_ sky130_fd_sc_hd__or3_1
X_10130_ net428 _05646_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] net749 _05572_ _05576_
+ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a2111oi_2
XANTENNA__09714__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16783__1327 vssd1 vssd1 vccd1 vccd1 _16783__1327/HI net1327 sky130_fd_sc_hd__conb_1
XFILLER_0_199_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13820_ net1150 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09469__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10963_ net379 _06474_ _06473_ net416 vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15224__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12702_ net365 net1877 net430 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__mux2_1
X_16470_ clknet_leaf_84_wb_clk_i net1588 _01278_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
X_13682_ _03199_ _03211_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__or2_1
X_10894_ _06110_ _06373_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15421_ clknet_leaf_12_wb_clk_i _01561_ _00229_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12633_ net1878 net345 net554 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__mux2_1
XANTENNA__12286__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10236__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15352_ clknet_leaf_77_wb_clk_i _01492_ _00165_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ net335 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\] net445 vssd1
+ vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_91_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11984__A0 _06626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14303_ net1108 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
X_11515_ team_02_WB.instance_to_wrap.top.pc\[6\] _06255_ team_02_WB.instance_to_wrap.top.pc\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_156_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15283_ clknet_leaf_68_wb_clk_i _01427_ _00096_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12495_ net320 net1716 net556 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09929__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14234_ net1095 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
X_11446_ net420 _06356_ _06516_ _06941_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__a31o_1
XANTENNA__11697__Y _07183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13103__A1_N net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14165_ net1242 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
X_11377_ _06872_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_189_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13116_ _07470_ _07514_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__and2_1
X_10328_ _05838_ _05840_ _05842_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__or4_1
X_14096_ net1226 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XANTENNA__10106__Y _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13047_ net790 _07332_ _07534_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__a211o_1
X_10259_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] net779 _05772_ _05773_
+ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14530__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08904__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1264 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__buf_2
XANTENNA__12969__B _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1251 net1252 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_2
Xfanout1262 net1263 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ net1135 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16737_ team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net177
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13949_ net1243 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16668_ clknet_leaf_66_wb_clk_i net1363 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.debounce_dly
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09880__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12196__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15619_ clknet_leaf_8_wb_clk_i _01759_ _00427_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_16599_ clknet_leaf_96_wb_clk_i _02718_ _01392_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10227__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09140_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\] net718 net688 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16715__1274 vssd1 vssd1 vccd1 vccd1 _16715__1274/HI net1274 sky130_fd_sc_hd__conb_1
XFILLER_0_161_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09632__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09071_ _04581_ _04587_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_20_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08022_ _03698_ _03702_ _03705_ _03701_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a22o_1
Xhold701 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11727__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold712 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold734 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold745 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _05442_ _04421_ net550 vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_139_Left_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10016__Y _05533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold789 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ net1047 _04215_ _04232_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a22o_1
XANTENNA__09699__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ net170 net1040 net1037 net1537 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout471_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A _07217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07806_ _03528_ _03484_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08786_ _04406_ _04409_ _04411_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__nor4_1
XFILLER_0_211_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07737_ _03424_ _03458_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout736_A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07668_ _03380_ _03382_ _03354_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_148_Left_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09871__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\] net678 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__a22o_1
X_07599_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout903_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09338_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] net929 net807 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\]
+ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a221o_1
XANTENNA__11415__C1 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09623__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\] net771 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a22o_1
X_11300_ net374 _06568_ _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12280_ net254 net1968 net570 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11162_ _06382_ _06638_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15219__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10941__B2 _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] net893 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a22o_1
X_11093_ _04951_ _06601_ _04950_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__a21oi_1
X_15970_ clknet_leaf_118_wb_clk_i _02110_ _00778_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12789__B _06398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14921_ net1216 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
X_10044_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\] net748 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__a22o_1
Xhold50 team_02_WB.instance_to_wrap.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 net1412
+ sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 _02583_ vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 team_02_WB.instance_to_wrap.ramstore\[17\] vssd1 vssd1 vccd1 vccd1 net1434
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1099 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
Xhold83 team_02_WB.instance_to_wrap.top.a1.data\[9\] vssd1 vssd1 vccd1 vccd1 net1445
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\] vssd1 vssd1 vccd1 vccd1
+ net1456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13803_ _03288_ net961 _03287_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__and3b_1
X_14783_ net1116 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11995_ net314 net2054 net480 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XANTENNA__11913__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16522_ clknet_leaf_0_wb_clk_i _02656_ _01329_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13734_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] _03242_ vssd1 vssd1 vccd1
+ vccd1 _03243_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10946_ _06270_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__or2_1
XANTENNA__10596__Y _06113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16453_ clknet_leaf_42_wb_clk_i net1408 _01261_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\]
+ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__and3_1
X_10877_ net373 _06077_ _06391_ net396 vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__o211a_1
XANTENNA__15751__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ net1981 net283 net553 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
X_15404_ clknet_leaf_2_wb_clk_i _01544_ _00212_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16384_ clknet_leaf_88_wb_clk_i _02519_ _01192_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13596_ net1464 net963 _03148_ net1067 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09614__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15335_ clknet_leaf_72_wb_clk_i _01478_ _00148_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12547_ net267 net2027 net444 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[25\]
+ _00079_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12478_ net252 net2151 net558 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ net1221 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13174__A2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ net794 _06924_ _06917_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15197_ net1246 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14148_ net1093 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XANTENNA__10932__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ net1108 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XANTENNA__14260__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_2
Xfanout1081 net1086 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_4
X_08640_ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_175_Right_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XANTENNA__15281__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08571_ team_02_WB.instance_to_wrap.top.a1.row1\[61\] _04237_ _04225_ vssd1 vssd1
+ vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11823__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09066__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09605__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ _04633_ _04635_ _04637_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_98_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08813__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12654__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16782__1326 vssd1 vssd1 vccd1 vccd1 _16782__1326/HI net1326 sky130_fd_sc_hd__conb_1
XFILLER_0_161_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] net758 net687 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08005_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03689_ _03721_ vssd1 vssd1
+ vccd1 vccd1 _03728_ sky130_fd_sc_hd__nand3_1
Xhold520 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold531 team_02_WB.instance_to_wrap.top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 net1893
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold542 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold564 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold575 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
X_09956_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\] net748 net710 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ net1486 _04435_ net930 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
X_09887_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\] net886 net858 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a22o_1
XANTENNA__11479__A2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1231 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ net157 net1042 net1034 net1407 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a22o_1
Xhold1242 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 team_02_WB.instance_to_wrap.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net2615
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1264 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1275 team_02_WB.instance_to_wrap.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net2637
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] net741 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ _04630_ net405 vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__nand2_1
X_11780_ net271 net2337 net595 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09844__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ _04349_ _04354_ _04344_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__and3b_1
XANTENNA__07855__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11034__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ _03044_ _03049_ _02768_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09057__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10662_ net996 _04421_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_123_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_62_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ net338 net2505 net458 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__mux2_1
XANTENNA__12564__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ net1469 net1013 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[10\]
+ sky130_fd_sc_hd__and2_1
X_10593_ _04462_ _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__nor2_4
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15120_ net1165 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
X_12332_ net327 net1712 net566 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10592__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15051_ net1233 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
X_12263_ net313 net2239 net574 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14002_ net1185 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
X_11214_ _06351_ _06718_ _06717_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_186_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11975__Y _07204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ net310 net2140 net577 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__mux2_1
XANTENNA__11908__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _06266_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11076_ _06574_ _06581_ _06582_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__or3_1
X_15953_ clknet_leaf_0_wb_clk_i _02093_ _00761_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_2
X_16714__1273 vssd1 vssd1 vccd1 vccd1 _16714__1273/HI net1273 sky130_fd_sc_hd__conb_1
X_10027_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] net831 net803 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\]
+ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__a221o_1
X_14904_ net1199 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
X_15884_ clknet_leaf_126_wb_clk_i _02024_ _00692_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10142__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14835_ net1073 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ net1082 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
X_11978_ net237 net2057 net478 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
XANTENNA__09296__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09835__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16505_ clknet_leaf_127_wb_clk_i _02639_ _01312_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929_ net371 _06326_ net398 vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__o21ai_1
X_13717_ _03204_ _03023_ net1066 _03200_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__and4b_1
X_14697_ net1214 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09048__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16436_ clknet_leaf_70_wb_clk_i net1538 _01244_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dfrtp_1
X_13648_ net1377 net1067 _03023_ _03194_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16367_ clknet_leaf_41_wb_clk_i _02507_ _01175_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13579_ team_02_WB.instance_to_wrap.top.a1.row1\[8\] _03110_ _03128_ team_02_WB.instance_to_wrap.top.a1.row1\[104\]
+ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15318_ clknet_leaf_72_wb_clk_i _01461_ _00131_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_16298_ clknet_leaf_37_wb_clk_i _02438_ _01106_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15249_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[8\]
+ _00062_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09220__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A1 _06134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] net929 net802 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a221o_1
XANTENNA__11818__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout307 _06891_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10905__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net320 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout329 _03568_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
X_09741_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\] net706 net700 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\]
+ _05254_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a221o_1
X_09672_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\] net810 net881 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10133__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08623_ net103 net1555 _04261_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
XANTENNA__12649__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _04217_ _04218_ net651 net793 net1680 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09287__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09826__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ _04179_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1176_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10964__Y _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12384__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09106_ _04613_ _04614_ _04615_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__or4_2
XFILLER_0_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\] net814 net895 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\]
+ _04548_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1131_X net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_211_Right_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold350 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold372 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10372__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 _04508_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_8
Xfanout841 _04403_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_4
Xfanout852 net854 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_8
X_09939_ _05449_ _05451_ _05453_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 _04543_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 _04539_ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_8
Xfanout885 _04537_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_4
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_4
X_12950_ team_02_WB.instance_to_wrap.top.pc\[15\] _06197_ vssd1 vssd1 vccd1 vccd1
+ _07470_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10124__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net360 net2406 net488 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
Xhold1061 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1083 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ _07398_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__or2_1
XANTENNA__12559__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1094 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13244__A _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ net344 net2428 net590 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
X_14620_ net1192 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XANTENNA__11690__C _07161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09278__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ net1186 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
X_11763_ net332 net1906 net597 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
XANTENNA__15232__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13502_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__or2_1
X_10714_ _06174_ _06230_ _06175_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__o21ai_1
X_14482_ net1177 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
X_11694_ _07130_ _07137_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__nand3_1
XFILLER_0_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13433_ _03040_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__inv_2
X_16221_ clknet_leaf_12_wb_clk_i _02361_ _01029_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__inv_2
XANTENNA__12294__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ clknet_leaf_121_wb_clk_i _02292_ _00960_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ net1943 net1018 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[26\]
+ sky130_fd_sc_hd__and2_1
X_10576_ _06090_ _06092_ net369 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__mux2_1
XANTENNA__09450__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ net259 net2267 net564 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__mux2_1
X_15103_ net1175 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16083_ clknet_leaf_57_wb_clk_i _02223_ _00891_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13295_ team_02_WB.instance_to_wrap.top.pc\[12\] net1053 _06908_ net935 vssd1 vssd1
+ vccd1 vccd1 _02997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ net1235 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12246_ net237 net2116 net575 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__mux2_1
XANTENNA__09202__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_75_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09175__Y _04692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ net642 _06278_ _06280_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_20_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_166_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11128_ _06353_ _06633_ _06632_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13301__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _06567_ _06568_ net412 vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15936_ clknet_leaf_110_wb_clk_i _02076_ _00744_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_16781__1325 vssd1 vssd1 vccd1 vccd1 _16781__1325/HI net1325 sky130_fd_sc_hd__conb_1
XANTENNA__10115__A2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ clknet_leaf_34_wb_clk_i _02007_ _00675_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12469__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11226__X _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13154__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14818_ net1191 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XANTENNA__13065__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09269__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15798_ clknet_leaf_21_wb_clk_i _01938_ _00606_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14749_ net1206 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12812__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12812__B2 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _03983_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_2__f_wb_clk_i_X clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16419_ clknet_leaf_80_wb_clk_i _02554_ _01227_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09441__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13540__A2 _03061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10354__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07985_ _03695_ net256 vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__and2b_1
X_09724_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\] net897 net941 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a22o_1
XANTENNA__10106__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\] net764 net707 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a22o_1
XANTENNA__12379__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ net90 net1523 net957 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09586_ net530 vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__inv_2
XFILLER_0_179_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08537_ _04171_ _04220_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout816_A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1179_X net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ net1580 net1006 net980 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1
+ vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08483__A1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09680__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire505 _05667_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_2
X_08399_ _04090_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__or3_1
Xwire516 _05439_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire527 _05146_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_2
X_10430_ _04997_ _05946_ _04993_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__a21oi_1
Xwire549 _04415_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_2
X_16713__1272 vssd1 vssd1 vccd1 vccd1 _16713__1272/HI net1272 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_150_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10361_ net390 _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__nor2_1
XANTENNA__15962__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ net1670 net337 net583 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
X_13080_ _07460_ _07524_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10292_ _05787_ _05807_ net968 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ net322 net1731 net474 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
Xhold180 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13239__A _02953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 team_02_WB.instance_to_wrap.ramaddr\[20\] vssd1 vssd1 vccd1 vccd1 net1553
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10345__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15227__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 net662 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_2
Xfanout671 _05964_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_2
XFILLER_0_205_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16770_ net1314 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_205_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout682 _04402_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_4
Xfanout693 _04394_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_70_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13982_ net1188 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XANTENNA__13295__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15721_ clknet_leaf_111_wb_clk_i _01861_ _00529_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12933_ team_02_WB.instance_to_wrap.top.pc\[26\] _06150_ vssd1 vssd1 vccd1 vccd1
+ _07453_ sky130_fd_sc_hd__nand2_1
XANTENNA__12289__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15652_ clknet_leaf_34_wb_clk_i _01792_ _00460_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13047__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ _05489_ _05491_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14603_ net1099 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
X_11815_ net280 net2243 net590 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
X_15583_ clknet_leaf_61_wb_clk_i _01723_ _00391_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12795_ _06102_ _07099_ _07317_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__and4_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11921__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ net264 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] net599 vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__mux2_1
X_14534_ net1213 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09671__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14465_ net1262 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
X_11677_ _05125_ _05978_ _07162_ _05973_ _05124_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ clknet_leaf_2_wb_clk_i _02344_ _01012_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13416_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] team_02_WB.instance_to_wrap.top.lcd.currentState\[0\]
+ _03023_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
X_10628_ team_02_WB.instance_to_wrap.top.pc\[27\] _06143_ vssd1 vssd1 vccd1 vccd1
+ _06145_ sky130_fd_sc_hd__and2_1
XANTENNA__09423__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14396_ net1192 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16135_ clknet_leaf_40_wb_clk_i _02275_ _00943_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08777__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13347_ net2635 net1015 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_106_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09974__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10559_ _04714_ net405 vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16066_ clknet_leaf_118_wb_clk_i _02206_ _00874_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13278_ net1635 net985 net967 _02988_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12229_ net2202 net305 net615 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__mux2_1
X_15017_ net1165 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_102_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13149__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10336__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07770_ _03451_ _03491_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__and3_1
X_15919_ clknet_leaf_44_wb_clk_i _02059_ _00727_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12199__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09440_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] net765 net693 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\]
+ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09371_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\] net921 net892 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_111_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _04015_ _04028_ _04032_ _04024_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_115_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07610__A team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08253_ _03967_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ _03892_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__B2 _04946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10019__Y _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12662__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1041_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout599_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1035_X net2397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _03648_ _03687_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__xor2_1
XANTENNA__10910__S net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\] net784 net712 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07899_ _03595_ _03619_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\] net919 net875 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] net781 net760 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11600_ net389 _07052_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11741__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12580_ net265 net1732 net440 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__mux2_1
XANTENNA__13208__A2_N net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09653__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ net419 _06635_ _06849_ net377 _07018_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__a221o_2
XFILLER_0_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14250_ net1117 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
X_11462_ _06007_ _06956_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09405__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13201_ net636 net936 net1020 net1400 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16780__1324 vssd1 vssd1 vccd1 vccd1 _16780__1324/HI net1324 sky130_fd_sc_hd__conb_1
XFILLER_0_190_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ _05927_ _05929_ _05420_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__o21a_1
XANTENNA__08759__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14181_ net1113 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
X_11393_ net1528 net307 net639 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XANTENNA__12572__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13132_ net229 _02897_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a21boi_1
X_10344_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\] net761 _05859_ _05860_
+ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a211o_1
XANTENNA_input62_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12144__Y _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _07529_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__xnor2_1
X_10275_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\] net832 net878 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a22o_1
XANTENNA__08070__B _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ net248 net2294 net476 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XANTENNA__09184__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11916__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__Y _04970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout490 _07196_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_8
X_16753_ net1297 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
X_13965_ net1248 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
X_15704_ clknet_leaf_121_wb_clk_i _01844_ _00512_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12916_ _04755_ _06147_ _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__a21o_1
X_16684_ clknet_leaf_65_wb_clk_i _02801_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09892__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ net1251 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
X_15635_ clknet_leaf_58_wb_clk_i _01775_ _00443_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ _05061_ _06186_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15566_ clknet_leaf_59_wb_clk_i _01706_ _00374_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _06720_ _06902_ _07299_ _07301_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and4_1
XFILLER_0_173_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14517_ net1257 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11729_ net330 net2393 net600 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
X_15497_ clknet_leaf_116_wb_clk_i _01637_ _00305_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15238__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14448_ net1232 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_211_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09947__A1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10791__A _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold905 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ net1125 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
Xhold916 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_2
Xhold927 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16118_ clknet_leaf_21_wb_clk_i _02258_ _00926_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap646 net647 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_2
Xhold949 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16049_ clknet_leaf_126_wb_clk_i _02189_ _00857_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_08940_ net1059 _04278_ _04315_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__or3b_2
XFILLER_0_177_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__A1 _06998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10309__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__A2 _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ net26 net1031 _04432_ net1623 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_209_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11826__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07822_ _03506_ _03541_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__xor2_2
XANTENNA__10190__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A _04588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _03457_ _03475_ _03460_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o21ai_1
X_16712__1271 vssd1 vssd1 vccd1 vccd1 _16712__1271/HI net1271 sky130_fd_sc_hd__conb_1
XFILLER_0_177_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07684_ _03363_ _03368_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__or2_1
X_09423_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\] net864 net855 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a221o_1
XANTENNA__12657__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14438__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_A _07187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__S net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13342__A net2352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09354_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\] net840 net675 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1089_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09635__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ _03976_ _03993_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10245__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16426__Q net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ net535 vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1256_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08236_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13195__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ _03879_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nor2_1
XANTENNA__12392__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ _03815_ _03816_ _03800_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout883_A _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_189_Right_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1152_X net2514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\] net760 net697 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_54_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11736__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10181__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Left_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ _06068_ _06094_ net394 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__mux2_1
X_13750_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03251_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12701_ net355 net1691 net432 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10893_ _05957_ net661 net658 _04653_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__a22o_1
X_13681_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\] _03198_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12567__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15420_ clknet_leaf_20_wb_clk_i _01560_ _00228_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_191_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12632_ net1665 net338 net555 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__mux2_1
XANTENNA__09626__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12563_ net328 net1833 net443 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__mux2_1
X_15351_ clknet_leaf_57_wb_clk_i _01491_ _00164_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15240__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _05604_ _06113_ _07006_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__o21ai_2
X_14302_ net1191 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12494_ net312 net1745 net556 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ clknet_leaf_70_wb_clk_i _01426_ _00095_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramaddr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11445_ net375 _06747_ _06940_ net382 vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_150_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15179__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14233_ net1096 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ net1193 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
X_11376_ net413 _06401_ _06853_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_189_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] net816 net804 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\]
+ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ team_02_WB.instance_to_wrap.top.pc\[16\] net1023 _02886_ net1028 vssd1 vssd1
+ vccd1 vccd1 _01497_ sky130_fd_sc_hd__a22o_1
X_14095_ net1226 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14811__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09157__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15680__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13046_ _07451_ _07533_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__and2_1
X_10258_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\] net840 net674 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a221o_1
Xfanout1230 net1236 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__buf_2
Xfanout1241 net1243 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_4
XFILLER_0_206_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10189_ _05699_ _05701_ _05703_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1252 net1255 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_2
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14997_ net1148 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
X_16736_ net1282 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13948_ net1243 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XANTENNA__09865__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16667_ clknet_leaf_66_wb_clk_i _00017_ _01409_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12477__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13879_ net1253 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15618_ clknet_leaf_101_wb_clk_i _01758_ _00426_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16598_ clknet_leaf_90_wb_clk_i _02717_ _01391_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15549_ clknet_leaf_13_wb_clk_i _01689_ _00357_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] net771 _04583_ _04585_
+ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08021_ _03733_ _03737_ _03742_ _03712_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a31o_2
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold702 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09396__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold713 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold724 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold746 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold768 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ net512 vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__inv_2
Xhold779 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14721__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09148__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] net959 vssd1 vssd1 vccd1
+ vccd1 _04444_ sky130_fd_sc_hd__or2_1
XANTENNA__08047__A2_N _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A _06865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net1467 net1039 net1037 team_02_WB.instance_to_wrap.ramstore\[10\] vssd1
+ vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1004_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10163__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ _03481_ _03494_ net366 vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_127_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\] net725 net673 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\]
+ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_197_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout464_A _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07736_ _03424_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _03388_ _03389_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__or2_1
XANTENNA__12387__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout729_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\] net739 net699 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\]
+ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07598_ team_02_WB.instance_to_wrap.top.a1.row2\[15\] net1010 _03321_ vssd1 vssd1
+ vccd1 vccd1 _02731_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09337_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] net823 net877 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_173_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\] net767 net746 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08219_ _03916_ _03918_ _03919_ _03926_ _03934_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o41ai_1
XANTENNA__16533__D net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09199_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\] net834 net903 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a22o_1
XANTENNA__11179__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ _06264_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _04993_ net661 net658 _04995_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14631__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09139__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] net899 net799 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\]
+ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a221o_1
X_11092_ _05976_ _06600_ _06022_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12789__C _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\] net753 net741 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a22o_1
X_14920_ net1112 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
XANTENNA__10223__X _05740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 net124 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__B2 net2352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold51 _02577_ vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_02_WB.instance_to_wrap.ramaddr\[8\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 _02579_ vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net1135 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15235__Q team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold84 net134 vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 net132 vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\]
+ _03284_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__and3_1
XFILLER_0_203_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14782_ net1128 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XANTENNA__09847__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ net304 net2617 net479 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XANTENNA__09311__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ clknet_leaf_5_wb_clk_i _02655_ _01328_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13733_ _03242_ net951 _03241_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_67_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12297__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ team_02_WB.instance_to_wrap.top.pc\[27\] _06269_ team_02_WB.instance_to_wrap.top.pc\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16452_ clknet_leaf_44_wb_clk_i net1389 _01260_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13664_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _03198_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_210_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10876_ net391 _06079_ _06080_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__or3_1
XFILLER_0_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15403_ clknet_leaf_15_wb_clk_i _01543_ _00211_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12615_ net1787 net270 net553 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
XANTENNA__11406__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16383_ clknet_leaf_88_wb_clk_i _02518_ _01191_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13595_ _03112_ _03135_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15334_ clknet_leaf_42_wb_clk_i _01477_ _00147_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12546_ net258 net2444 net442 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15265_ clknet_leaf_80_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[24\]
+ _00078_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12477_ net238 net2460 net556 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16711__1270 vssd1 vssd1 vccd1 vccd1 _16711__1270/HI net1270 sky130_fd_sc_hd__conb_1
XANTENNA_4 _04371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09378__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14216_ net1113 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
X_11428_ net420 _06481_ _06922_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a21o_1
X_15196_ net1246 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14147_ net1136 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
X_11359_ _06201_ _06206_ _06208_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_169_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ net1127 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13029_ _07352_ _07440_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_206_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10145__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15426__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 team_02_WB.instance_to_wrap.top.a1.instruction\[12\] vssd1 vssd1 vccd1
+ vccd1 net1060 sky130_fd_sc_hd__buf_2
Xfanout1071 net61 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_2
XANTENNA__09550__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1085 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_4
Xfanout1093 net1094 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_2
XFILLER_0_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08570_ net1010 _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11645__B1 _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16719_ net1351 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09302__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12000__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09122_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\] net808 net902 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\]
+ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12507__Y _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] net755 net731 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08004_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03689_ _03721_ vssd1 vssd1
+ vccd1 vccd1 _03727_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold521 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold532 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold543 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12670__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\] net756 net680 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout581_A _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net1047 _04190_ _04202_ net1009 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__a32o_1
XANTENNA__10136__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\] net918 net862 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a22o_1
Xhold1210 team_02_WB.instance_to_wrap.ramload\[3\] vssd1 vssd1 vccd1 vccd1 net2572
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1232 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net158 net1040 net1037 net1514 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
Xhold1254 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1265 team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1 net2627
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net2638
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1115_X net2477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08768_ net846 _04365_ _04370_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and3_4
XFILLER_0_197_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07719_ _03440_ _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__nor2_1
X_08699_ _04276_ _04320_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10730_ net994 net848 vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10661_ team_02_WB.instance_to_wrap.top.pc\[22\] _06177_ vssd1 vssd1 vccd1 vccd1
+ _06178_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ net332 net1819 net458 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13380_ net2638 net1014 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.next_FetchedData\[9\]
+ sky130_fd_sc_hd__and2_1
X_10592_ _04463_ _04467_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12331_ net321 net2525 net564 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11050__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15050_ net1235 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_12262_ net304 net2160 net573 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ net409 _06480_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__nand2_1
X_14001_ net1231 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_186_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12193_ net302 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] net579 vssd1
+ vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12580__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ team_02_WB.instance_to_wrap.top.pc\[21\] _06265_ team_02_WB.instance_to_wrap.top.pc\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09780__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11075_ _04865_ _06026_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__xnor2_1
X_15952_ clknet_leaf_23_wb_clk_i _02092_ _00760_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10127__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\] net904 net872 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a22o_1
X_14903_ net1210 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XANTENNA__09532__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ clknet_leaf_114_wb_clk_i _02023_ _00691_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11924__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15192__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14834_ net1177 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14765_ net1121 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
X_11977_ net246 net1478 net479 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16504_ clknet_leaf_1_wb_clk_i _02638_ _01311_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13716_ net1585 _03231_ _03232_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__o21a_1
X_10928_ net391 _06315_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14696_ net1111 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16435_ clknet_leaf_64_wb_clk_i _02570_ _01243_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09048__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ _03289_ _03114_ _03115_ _03193_ _03023_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a311oi_1
X_10859_ _04693_ _05956_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09599__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16366_ clknet_leaf_46_wb_clk_i _02506_ _01174_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_167_Left_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ team_02_WB.instance_to_wrap.top.a1.row1\[56\] _03117_ _03119_ team_02_WB.instance_to_wrap.top.a1.row1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15317_ clknet_leaf_70_wb_clk_i _01460_ _00130_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramstore\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10602__B2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ net324 net1647 net446 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
XANTENNA__16224__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16297_ clknet_leaf_112_wb_clk_i _02437_ _01105_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08079__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15248_ clknet_leaf_104_wb_clk_i team_02_WB.instance_to_wrap.top.ru.next_FetchedInstr\[7\]
+ _00061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12490__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15179_ net1145 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XANTENNA__10366__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10905__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15204__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire647_A _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_0_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09740_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\] net754 net727 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a22o_1
XANTENNA__10118__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

