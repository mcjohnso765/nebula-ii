* NGSPICE file created from team_01_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt team_01_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10669__A1 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] net848
+ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and3_1
XANTENNA__08731__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\] net629 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\]
+ _04884_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08709__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08553_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] net748 net715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\]
+ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a221o_1
XANTENNA__13083__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08484_ net1108 net1111 net1114 net1106 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12665__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1071_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A _08024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09105_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\] net752 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\]
+ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1336_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09036_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] net729 net718 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15277__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold340 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\] vssd1 vssd1 vccd1 vccd1
+ net1956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 net83 vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12897__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold373 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09706__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 _03321_ vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net821 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
XANTENNA__08970__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 net832 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_4
X_09938_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\] net914 vssd1
+ vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__and3_1
Xfanout842 net844 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout853 _04760_ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout864 net866 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_2
Xfanout886 net889 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
Xfanout897 net900 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__clkbuf_2
X_09869_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\] net693 _06115_ _06117_
+ _06118_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1040 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11900_ net494 _07846_ _08008_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12880_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] vssd1 vssd1 vccd1
+ vccd1 _03589_ sky130_fd_sc_hd__or2_2
Xhold1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1084 _02070_ vssd1 vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13244__B net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ net2603 net249 net480 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14550_ net1332 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11762_ net781 _07896_ _07895_ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_83_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13501_ _03846_ _03848_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ net521 _06976_ _06971_ _06969_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__o211a_1
X_14481_ net1380 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
XANTENNA__12575__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ team_01_WB.instance_to_wrap.cpu.K0.count\[0\] team_01_WB.instance_to_wrap.cpu.K0.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__nand2b_1
XANTENNA__14356__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16220_ clknet_leaf_42_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[1\]
+ _00088_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13432_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _06415_ vssd1 vssd1 vccd1
+ vccd1 _03785_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10644_ _06907_ _06901_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18201__1575 vssd1 vssd1 vccd1 vccd1 _18201__1575/HI net1575 sky130_fd_sc_hd__conb_1
XANTENNA__08789__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16151_ net1322 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10575_ _04907_ _04957_ _04906_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__o21ba_1
X_13363_ net2 net800 net595 net2932 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15102_ net1293 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16397__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12314_ net1955 net250 net429 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__mux2_1
X_16082_ net1405 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13294_ net131 net810 net805 net1717 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17642__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11919__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13534__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ net1190 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ net2005 net284 net435 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09753__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ net3032 net198 net443 vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08961__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _07388_ _07390_ net541 vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__mux2_1
XANTENNA__17792__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10124__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16984_ clknet_leaf_29_wb_clk_i _02544_ _00847_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_15935_ net1340 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__inv_2
X_11058_ _07075_ _07311_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_60_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10009_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\] net722 _06251_ _06253_
+ _06255_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13435__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15866_ net1307 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__inv_2
XANTENNA__17022__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17605_ clknet_leaf_135_wb_clk_i _03165_ _01468_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14817_ net1352 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13065__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15797_ net1173 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__inv_2
XANTENNA__14262__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17536_ clknet_leaf_140_wb_clk_i _03096_ _01399_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14748_ net1273 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13470__C1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10823__A1 _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17467_ clknet_leaf_37_wb_clk_i _03027_ _01330_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12485__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14679_ net1364 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XANTENNA__17172__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16418_ clknet_leaf_102_wb_clk_i net2841 _00281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17398_ clknet_leaf_30_wb_clk_i _02958_ _01261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ clknet_leaf_66_wb_clk_i net1854 _00217_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10051__A2 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18019_ net1596 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XANTENNA__11829__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09095__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13329__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09526__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08430__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\] _04661_ _05964_
+ _05969_ _05970_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09823__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout377_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09654_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\] net744 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08605_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] net730 _04857_
+ _04858_ _04865_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09585_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] net753 net695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\]
+ _05835_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a221o_1
XANTENNA__09261__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout544_A _06315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08536_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\] net961
+ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10200__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12395__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net1106 net1108 net1111 net1114 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout711_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout809_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08398_ net1118 net943 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__and2_4
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13764__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14904__A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10042__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\] net942 vssd1
+ vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09019_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\] net953 vssd1
+ vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__and3_1
X_10291_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] net859 vssd1
+ vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12030_ net2624 net309 net466 vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold170 net94 vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold181 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1 vccd1 net1797
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09436__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 net96 vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09733__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout661 _04737_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_8
Xfanout672 _04729_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13981_ _04169_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__inv_2
Xfanout683 _04696_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_6
Xfanout694 _04690_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_6
X_15720_ net1208 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
X_12932_ net364 _03625_ _03626_ net1053 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__a32o_1
XANTENNA__10502__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15651_ net1220 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
X_12863_ net1156 team_01_WB.instance_to_wrap.cpu.DM0.enable team_01_WB.instance_to_wrap.cpu.DM0.state\[0\]
+ net766 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__or4bb_1
XANTENNA__13047__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14244__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14602_ net1411 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
X_11814_ net2519 net280 net480 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15582_ net1291 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
X_12794_ net2436 net210 net378 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
X_17321_ clknet_leaf_42_wb_clk_i _02881_ _01184_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14533_ net1320 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11745_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] net674 net774 vssd1 vssd1
+ vccd1 vccd1 _07883_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17252_ clknet_leaf_128_wb_clk_i _02812_ _01115_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14464_ net1390 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11676_ net2044 net1159 vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ clknet_leaf_95_wb_clk_i _01870_ _00071_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_13415_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _06827_ vssd1 vssd1
+ vccd1 vccd1 _03768_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10627_ _06108_ _06071_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__and2b_1
X_17183_ clknet_leaf_0_wb_clk_i _02743_ _01046_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08226__A2 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14395_ net1352 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16134_ net1314 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11230__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ net10 net801 net596 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1
+ vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a22o_1
X_10558_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\] net626 net622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\]
+ _06821_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08812__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16065_ net1368 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__inv_2
X_13277_ net80 net810 net597 net1734 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10489_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] net847
+ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13936__A_N net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15016_ net1181 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
X_12228_ net3214 net311 net442 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12159_ net1922 net243 net449 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
XANTENNA__10741__A0 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09643__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13286__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16967_ clknet_leaf_126_wb_clk_i _02527_ _00830_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_15918_ net1380 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__inv_2
X_16898_ clknet_leaf_144_wb_clk_i _02458_ _00761_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08162__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15849_ net1221 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_133_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13038__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09370_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] net956 vssd1
+ vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10020__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16562__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08321_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\] net3113 net1051 vssd1 vssd1
+ vccd1 vccd1 _03426_ sky130_fd_sc_hd__mux2_1
X_17519_ clknet_leaf_93_wb_clk_i _03079_ _01382_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13104__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08252_ net2399 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\] net1046 vssd1 vssd1
+ vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08425__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _04580_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10029__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09818__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11772__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17068__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14171__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09256__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout759_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] net957
+ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and3_1
X_18200__1574 vssd1 vssd1 vccd1 vccd1 _18200__1574/HI net1574 sky130_fd_sc_hd__conb_1
XFILLER_0_39_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08153__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16905__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] net942
+ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13029__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] net917 vssd1
+ vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08519_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] net653 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\]
+ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a221o_1
XANTENNA__10799__A0 _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\] net924 vssd1
+ vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and3_1
XANTENNA__13014__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07765_ vssd1 vssd1 vccd1 vccd1
+ _07767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11461_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] net1063 _07711_ vssd1 vssd1 vccd1
+ vccd1 _07714_ sky130_fd_sc_hd__and3_1
XANTENNA__12853__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ net1646 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\] net826 vssd1 vssd1
+ vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10412_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] net913 vssd1
+ vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__and3_1
XANTENNA__11212__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ _04332_ _04334_ _04336_ _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__or4_1
X_11392_ _07243_ _07265_ _07568_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12960__A1 _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ net2947 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\] net824 vssd1 vssd1
+ vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
XANTENNA__12960__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ _06037_ _06605_ _05488_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10971__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09169__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14162__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\] net630 _06535_ _06536_
+ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__a2111o_1
X_13062_ net1751 net834 net354 _03694_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XANTENNA_input55_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net2373 net283 net463 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
XANTENNA__16435__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1401 net1402 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__buf_4
X_17870_ clknet_leaf_96_wb_clk_i _03420_ _01690_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1412 net1413 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10105__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09463__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16821_ clknet_leaf_8_wb_clk_i _02381_ _00684_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13268__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 net482 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout491 _08025_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_4
X_16752_ clknet_leaf_25_wb_clk_i _02312_ _00615_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13964_ _04148_ _04154_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15703_ net1247 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
X_12915_ net2109 net604 net586 _03614_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
X_16683_ clknet_leaf_56_wb_clk_i _02243_ _00546_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10121__B _06382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ net3266 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[8\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_88_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11932__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15634_ net1184 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
X_12846_ net2312 net275 net368 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08807__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ net1213 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
XANTENNA__13432__B _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08447__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ net2016 net250 net377 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17304_ clknet_leaf_28_wb_clk_i _02864_ _01167_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ net1403 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17980__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10254__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11728_ _07867_ _07868_ net777 vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15496_ net1181 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17235_ clknet_leaf_49_wb_clk_i _02795_ _01098_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ net1385 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11659_ net2577 net1158 net569 net1113 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__a22o_1
XANTENNA__12763__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18016__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__C1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10006__A2 _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__B _07456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17166_ clknet_leaf_53_wb_clk_i _02726_ _01029_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14378_ net1382 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08542__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold906 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold917 team_01_WB.instance_to_wrap.cpu.f0.num\[24\] vssd1 vssd1 vccd1 vccd1 net2533
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__A1 team_01_WB.instance_to_wrap.a1.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16117_ net1364 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__inv_2
Xhold928 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _03746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17097_ clknet_leaf_40_wb_clk_i _02657_ _00960_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold939 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14153__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16048_ net1377 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17360__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ net1116 net763 net590 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a21o_1
Xhold1606 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1617 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16928__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1628 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\] vssd1 vssd1 vccd1 vccd1
+ net3244 sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ clknet_leaf_62_wb_clk_i _03548_ _01819_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1639 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3255 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11408__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12003__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12938__S net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14208__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09422_ _05652_ _05685_ net582 vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__mux2_2
XANTENNA__10493__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09353_ _05608_ _05614_ _05615_ _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08438__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__mux2_1
XANTENNA__10245__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09284_ _05539_ _05540_ _05546_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08235_ net1821 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12673__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ net1740 net550 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1
+ vccd1 vccd1 _03529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11745__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16458__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08097_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] _04488_ team_01_WB.instance_to_wrap.cpu.f0.num\[6\]
+ _04479_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold1357_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14144__B1 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08999_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] net857 vssd1
+ vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__and3_1
XANTENNA__09714__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17853__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13009__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10222__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10961_ _05487_ _06606_ _06608_ _05348_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__o211ai_1
XANTENNA__08677__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12848__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13533__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net2219 net240 net385 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__mux2_1
XANTENNA__09730__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ net772 _07464_ _07477_ net968 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a31o_1
XANTENNA__10484__A2 _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10892_ _05206_ _07155_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12631_ net2414 net196 net393 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ net1303 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ net2416 net290 net404 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17233__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ net1908 _04444_ net1172 vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__o21ai_1
X_11513_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] _07754_ _07755_ vssd1 vssd1 vccd1
+ vccd1 _03369_ sky130_fd_sc_hd__a21bo_1
X_15281_ net1195 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XANTENNA__12583__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ net2452 net313 net414 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
X_17020_ clknet_leaf_13_wb_clk_i _02580_ _00883_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09458__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14232_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\] _04250_ _04278_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\]
+ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11444_ _07697_ net3259 _07685_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12933__B2 _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\] _04256_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\]
+ _04312_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__a221o_1
X_11375_ _07004_ _07330_ _07638_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14135__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] net1161 vssd1 vssd1 vccd1 vccd1
+ _03727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10326_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] net709 net757 vssd1
+ vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14094_ net790 net788 _04241_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__and3_4
XFILLER_0_46_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11927__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17922_ clknet_leaf_78_wb_clk_i net3095 _01742_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\]
+ sky130_fd_sc_hd__dfrtp_1
X_13045_ _06826_ net571 net358 vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10257_ net582 _06486_ _06487_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1220 net1227 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09193__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1231 net1235 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10188_ net579 _06450_ _06416_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13427__B _06348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1242 net1245 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
X_17853_ clknet_leaf_104_wb_clk_i _03403_ _01673_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1253 net1268 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1264 net1268 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_2
Xfanout1275 net1276 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_2
X_16804_ clknet_leaf_129_wb_clk_i _02364_ _00667_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10132__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1286 net1289 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__buf_4
Xfanout1297 net1300 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__buf_4
XANTENNA__13646__C1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17784_ clknet_leaf_113_wb_clk_i _03342_ _01605_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14996_ net1238 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XANTENNA__08117__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13110__A1 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13947_ net1164 net1057 net3267 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[28\]
+ sky130_fd_sc_hd__and3b_1
X_16735_ clknet_leaf_2_wb_clk_i _02295_ _00598_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12758__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10475__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16666_ clknet_leaf_106_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[20\]
+ _00529_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11672__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13878_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__inv_2
XANTENNA__08537__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15617_ net1289 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
X_12829_ net2586 net195 net367 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16597_ clknet_leaf_57_wb_clk_i _02225_ _00460_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ net1235 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12493__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15479_ net1243 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17218_ clknet_leaf_0_wb_clk_i _02778_ _01081_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09368__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18198_ net1572 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
XFILLER_0_13_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12924__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08703__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17149_ clknet_leaf_127_wb_clk_i _02709_ _01012_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold714 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\] vssd1 vssd1 vccd1 vccd1
+ net2330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10307__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold725 team_01_WB.instance_to_wrap.cpu.f0.num\[23\] vssd1 vssd1 vccd1 vccd1 net2341
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\] vssd1 vssd1 vccd1 vccd1
+ net2352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] _04777_ _06218_
+ _06221_ _06225_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a2111o_1
Xhold769 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17876__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] net884 vssd1
+ vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__and3_1
XANTENNA__13618__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08853_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\] net907 vssd1
+ vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09534__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1403 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3019 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout192_A _07874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1414 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net3030
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17106__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1425 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1436 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\] vssd1 vssd1 vccd1 vccd1
+ net3052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08784_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] net856
+ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and3_1
Xhold1458 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3074 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08108__A1 _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1469 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3085 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08108__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13101__B2 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12668__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout457_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11663__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09405_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\] net896 vssd1
+ vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1366_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10218__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] net878
+ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09267_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\] net891 vssd1
+ vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__and3_1
XANTENNA__16280__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14184__A _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08831__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08218_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] net845
+ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and3_1
XANTENNA__09709__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12915__B2 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08149_ net1811 net551 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1
+ vccd1 vccd1 _03546_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14912__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09792__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _06319_ _06597_ _06869_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08910__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] net608 _06358_ _06360_
+ _06362_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_105_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11091_ _06109_ _07354_ _07020_ _06971_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13528__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] net630 _06280_ _06296_
+ _06299_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09544__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold30 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\] vssd1 vssd1 vccd1 vccd1 net1646
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] vssd1 vssd1 vccd1 vccd1 net1657
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 net1668
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1350 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold63 team_01_WB.instance_to_wrap.cpu.DM0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1679
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold74 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\] vssd1 vssd1 vccd1 vccd1
+ net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 net1701
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold96 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[18\] vssd1 vssd1 vccd1 vccd1 net1712
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09741__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13801_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] team_01_WB.instance_to_wrap.cpu.f0.i\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14781_ net1396 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
XANTENNA__12578__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net2770 net244 net468 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13643__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ clknet_leaf_73_wb_clk_i _02148_ _00383_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13732_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _04018_ vssd1 vssd1 vccd1 vccd1
+ _04049_ sky130_fd_sc_hd__or2_1
X_10944_ _07206_ _07207_ net528 vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11654__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16451_ clknet_leaf_101_wb_clk_i _02079_ _00314_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_13663_ _07981_ _03990_ net188 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10875_ net523 _07041_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__nand2_2
XFILLER_0_116_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17749__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15402_ net1198 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XANTENNA__10209__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12614_ net2014 net215 net395 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
X_16382_ clknet_leaf_115_wb_clk_i net1163 _00250_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09075__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net768 _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_85_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18121_ net1495 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15333_ net1226 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
X_12545_ net1871 net254 net404 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08822__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13202__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09188__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18052_ net1614 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15264_ net1287 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XANTENNA__08092__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12476_ net2793 net224 net413 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17003_ clknet_leaf_60_wb_clk_i _02563_ _00866_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17899__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14215_ net2104 net584 _04372_ net1170 vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__o211a_1
X_11427_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\] net1162 _04577_ _07683_ vssd1
+ vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__a22o_1
XANTENNA_5 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15195_ net1318 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10127__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08586__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14108__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__A3 _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _04158_ _04305_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11358_ _07620_ _07621_ _07615_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__and3b_1
XFILLER_0_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17129__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] net946 vssd1
+ vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__and3_1
X_14077_ net793 _04226_ net787 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__and3_4
XFILLER_0_123_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11289_ _07010_ _07014_ net529 vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__mux2_1
XANTENNA__12874__B1_N net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13028_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\] _03671_ net1029 vssd1
+ vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__mux2_1
X_17905_ clknet_leaf_107_wb_clk_i _03455_ _01725_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_wire258_A _07929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 net1052 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
X_18079__1453 vssd1 vssd1 vccd1 vccd1 _18079__1453/HI net1453 sky130_fd_sc_hd__conb_1
Xfanout1061 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 net1061
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11893__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17836_ clknet_leaf_87_wb_clk_i net837 _01657_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1072 net1076 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_2
Xfanout1083 net1085 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17279__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12488__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17767_ clknet_leaf_97_wb_clk_i _03325_ _01588_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14979_ net1219 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
X_16718_ clknet_leaf_50_wb_clk_i _02278_ _00581_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10448__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17698_ clknet_leaf_71_wb_clk_i _03258_ _01537_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11197__A1_N _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16649_ clknet_leaf_87_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[3\]
+ _00512_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13901__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] net893
+ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__and3_1
XANTENNA__13112__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09052_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\] net856
+ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09529__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08433__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] vssd1 vssd1 vccd1 vccd1
+ net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold533 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\] vssd1 vssd1 vccd1 vccd1
+ net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13570__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09826__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold577 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] net893 vssd1
+ vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__and3_1
Xhold599 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1114_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08905_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] net852 vssd1
+ vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__and3_1
X_09885_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] net870 vssd1
+ vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__and3_1
XANTENNA__09264__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1200 team_01_WB.instance_to_wrap.cpu.K0.code\[6\] vssd1 vssd1 vccd1 vccd1 net2816
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\] vssd1 vssd1 vccd1 vccd1
+ net2827 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13782__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1222 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\] net850
+ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1233 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10203__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1255 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09561__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1266 team_01_WB.instance_to_wrap.a1.ADR_I\[24\] vssd1 vssd1 vccd1 vccd1 net2882
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12398__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1277 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\] net753 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\]
+ _05019_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a221o_1
Xhold1288 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\] vssd1 vssd1 vccd1 vccd1
+ net2904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10439__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08698_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\] net935
+ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13389__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10660_ _05345_ _05309_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08905__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] net760 _05581_ _05582_
+ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a22o_4
XFILLER_0_10_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ net1156 net765 _06850_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 _06854_
+ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12330_ net2193 net292 net430 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12261_ net3224 net312 net438 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15738__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__C1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _04184_ _04185_ _04172_ _04180_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a2bb2o_1
X_11212_ net538 _07475_ _07471_ _06996_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__a211o_1
XANTENNA__09736__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08640__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ net2310 net243 net445 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11143_ _05448_ _05515_ _05583_ net548 net503 net518 vssd1 vssd1 vccd1 vccd1 _07407_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__09517__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_132_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_15951_ net1391 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__inv_2
XANTENNA__17421__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11074_ net321 _07330_ _07337_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10025_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\] net908 vssd1
+ vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and3_1
X_14902_ net1306 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15882_ net1356 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09471__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17621_ clknet_leaf_26_wb_clk_i _03181_ _01484_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10912__A1_N net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ net1339 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13616__A2 _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11506__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17552_ clknet_leaf_23_wb_clk_i _03112_ _01415_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14764_ net1257 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XANTENNA__08087__A team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10410__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ net3044 net287 net467 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16503_ clknet_leaf_75_wb_clk_i net3049 _00366_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_13715_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] _04035_ net783 vssd1 vssd1
+ vccd1 vccd1 _01852_ sky130_fd_sc_hd__mux2_1
X_17483_ clknet_leaf_46_wb_clk_i _03043_ _01346_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ _05205_ net342 _07184_ _07185_ _07176_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14695_ net1372 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11940__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13721__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13646_ net187 _03976_ _03977_ net772 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16434_ clknet_leaf_107_wb_clk_i _02062_ _00297_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ _06607_ _06612_ _06833_ _05212_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10850__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16365_ clknet_leaf_65_wb_clk_i net1770 _00233_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
X_13577_ _03841_ _03850_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__nor2_1
X_10789_ _07051_ _07052_ net515 vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15316_ net1237 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
X_18104_ net1478 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
X_12528_ net2071 net295 net410 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__mux2_1
X_16296_ clknet_leaf_111_wb_clk_i _01930_ _00164_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ net1601 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
X_15247_ net1248 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XANTENNA__15648__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ net2724 net260 net417 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
XANTENNA__12771__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16519__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11895__B _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ net1198 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14129_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\] _04238_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\]
+ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__a22o_1
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10118__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09670_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\] net898 vssd1
+ vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17914__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10023__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\] _04753_ net619
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] vssd1 vssd1 vccd1 vccd1
+ _04885_ sky130_fd_sc_hd__a22o_1
X_17819_ clknet_leaf_66_wb_clk_i _03376_ _01640_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] net721 net701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12011__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08428__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ net1084 net878 vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14727__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09039__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout322_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1064_A team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] net916 vssd1
+ vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09259__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09035_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] net751 net721 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\]
+ _05286_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12681__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1231_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1329_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16199__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold330 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _02104_ vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17444__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08460__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 _02000_ vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold385 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__buf_2
Xfanout821 net833 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_2
Xfanout832 net833 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_2
X_09937_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\] net958 vssd1
+ vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__and3_1
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_4
XANTENNA__13806__A team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09868_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] net753 _06112_ _06120_
+ _06122_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__a2111o_1
Xfanout887 _04742_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_4
Xhold1030 team_01_WB.instance_to_wrap.cpu.K0.code\[7\] vssd1 vssd1 vccd1 vccd1 net2646
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net902 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_4
Xhold1041 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09291__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1052 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\] net945 vssd1
+ vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__and3_1
XANTENNA__13059__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1063 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] vssd1 vssd1 vccd1 vccd1
+ net2679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _06059_ _06060_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or4_1
Xhold1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13017__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1096 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net780 _07952_ _07951_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__a21o_4
XANTENNA__09278__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14271__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11045__B _06933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11761_ _04483_ _07653_ net674 vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__mux2_1
XANTENNA__12856__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _05134_ _05167_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a22o_1
X_10712_ _06973_ _06975_ net515 vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14480_ net1380 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
X_11692_ net3012 net155 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13431_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _06526_ _07672_ _07671_
+ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10643_ _05757_ _06905_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16150_ net1332 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__inv_2
X_18078__1452 vssd1 vssd1 vccd1 vccd1 _18078__1452/HI net1452 sky130_fd_sc_hd__conb_1
X_13362_ net13 net802 _03747_ net2370 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
X_10574_ _06615_ _06778_ _06834_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__a31o_1
XANTENNA__09450__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15101_ net1281 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ net2544 net257 net428 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12591__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16081_ net1376 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13293_ net132 net811 net805 net1738 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13534__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15032_ net1259 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
X_12244_ net2930 net224 net436 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__mux2_1
XANTENNA__09466__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__A _04624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ net3146 net286 net443 vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16811__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10405__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17937__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11126_ _07231_ _07389_ net522 vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16983_ clknet_leaf_9_wb_clk_i _02543_ _00846_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11935__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13716__A team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15934_ net1342 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__inv_2
X_11057_ _07105_ _07320_ net534 vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10008_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\] net703 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13435__B _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09632__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15865_ net1193 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17604_ clknet_leaf_138_wb_clk_i _03164_ _01467_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14816_ net1357 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
X_15796_ net1237 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14262__A2 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17535_ clknet_leaf_4_wb_clk_i _03095_ _01398_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14747_ net1295 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
X_11959_ net2736 net301 net473 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XANTENNA__12766__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10284__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13451__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17466_ clknet_leaf_36_wb_clk_i _03026_ _01329_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10823__A2 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14678_ net1378 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XANTENNA__08545__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16417_ clknet_leaf_98_wb_clk_i _02045_ _00280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\]
+ sky130_fd_sc_hd__dfstp_1
X_13629_ net969 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _03962_ _03963_
+ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
X_17397_ clknet_leaf_9_wb_clk_i _02957_ _01260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09977__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16348_ clknet_leaf_65_wb_clk_i net1739 _00216_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XANTENNA__17467__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10587__A1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09441__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15378__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ clknet_leaf_71_wb_clk_i _01916_ _00147_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10018__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09729__B1 _05991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18018_ net1595 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16491__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12006__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09722_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] net738 net692 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a22o_1
X_09653_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\] net722 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a22o_1
XANTENNA__09542__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_A _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\] net740 net703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a22o_1
XANTENNA__15841__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ _05834_ _05845_ _05846_ _05847_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or4_1
XANTENNA__14253__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ _04797_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12676__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11067__A2 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout537_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1279_A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ net1017 net911 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nand2_1
XANTENNA__08455__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08397_ net971 net948 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and2_4
XANTENNA_fanout704_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09968__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__C1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18033__1599 vssd1 vssd1 vccd1 vccd1 net1599 _18033__1599/LO sky130_fd_sc_hd__conb_1
XANTENNA__11775__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10924__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] net928
+ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10290_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\] net895 vssd1
+ vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold160 _02002_ vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _02010_ vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\] vssd1 vssd1 vccd1 vccd1
+ net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold193 _02012_ vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout640 _04757_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_8
Xfanout651 _04747_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_6
XANTENNA__13536__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_8
X_13980_ net1170 _04168_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__nand2_2
Xfanout673 _04729_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
Xfanout684 _04696_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout695 _04688_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_6
X_12931_ net1026 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] vssd1 vssd1 vccd1
+ vccd1 _03626_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13970__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12862_ team_01_WB.instance_to_wrap.a1.WRITE_I team_01_WB.instance_to_wrap.cpu.RU0.state\[1\]
+ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__or3_2
X_15650_ net1289 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14244__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14601_ net1404 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ net776 _07936_ _07937_ _07938_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_69_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15581_ net1282 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
X_12793_ net2124 net291 net376 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XANTENNA__12586__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13452__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14532_ net1323 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
X_17320_ clknet_leaf_45_wb_clk_i _02880_ _01183_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11744_ net675 _07640_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08365__A team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ net1390 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XANTENNA__12007__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17251_ clknet_leaf_133_wb_clk_i _02811_ _01114_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11675_ net1709 net1159 vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13414_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _06827_ vssd1 vssd1
+ vccd1 vccd1 _03767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16202_ clknet_leaf_95_wb_clk_i _01869_ _00070_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _06600_ _06889_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__and2_1
X_17182_ clknet_leaf_3_wb_clk_i _02742_ _01045_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14394_ net1380 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ net1320 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ net11 net801 net596 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1
+ vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08631__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\] net650 net633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13210__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09196__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ net1374 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__inv_2
X_13276_ net81 net810 net597 net1849 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] net759 _06750_ _06751_
+ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__a22o_2
X_15015_ net1180 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
X_12227_ net2422 net261 net441 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XANTENNA__10135__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09924__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ net2440 net316 net447 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XANTENNA__10741__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _05889_ net335 net331 _06039_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__o2bb2a_1
X_12089_ net2047 net264 net456 vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
X_16966_ clknet_leaf_140_wb_clk_i _02526_ _00829_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_15917_ net1381 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__inv_2
XANTENNA__09362__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16897_ clknet_leaf_136_wb_clk_i _02457_ _00760_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15848_ net1219 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__inv_2
XANTENNA__10301__C _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12496__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15779_ net1219 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XANTENNA__13443__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17518_ clknet_leaf_55_wb_clk_i _03078_ _01381_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_08251_ net2859 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
XANTENNA__08706__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17449_ clknet_leaf_42_wb_clk_i _03009_ _01312_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16857__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13746__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _04564_ _04571_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08622__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13120__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09537__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1027_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16237__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09705_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] net962 vssd1
+ vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__and3_1
XANTENNA__09272__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18077__1451 vssd1 vssd1 vccd1 vccd1 _18077__1451/HI net1451 sky130_fd_sc_hd__conb_1
XANTENNA_fanout654_A _04743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1396_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09636_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\] net941 vssd1
+ vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__and3_1
XANTENNA__15571__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14226__A2 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17632__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ net1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] net955 vssd1
+ vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10919__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08518_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\] net627 net611 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09498_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] net941 vssd1
+ vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18215__1586 vssd1 vssd1 vccd1 vccd1 _18215__1586/HI net1586 sky130_fd_sc_hd__conb_1
XFILLER_0_37_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09653__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__A1 _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08449_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17782__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ net1063 _07711_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08913__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\] net956 vssd1
+ vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11391_ _07197_ _07307_ _07625_ _07640_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ net2528 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] net819 vssd1 vssd1
+ vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
X_10342_ _06037_ _06605_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13061_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\] _03693_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__mux2_1
XANTENNA__15746__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10273_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] net884 vssd1
+ vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and3_1
XANTENNA__14650__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12012_ net2043 net222 net465 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
XANTENNA__09744__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1402 net1413 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__buf_4
Xfanout1413 net1414 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17162__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16820_ clknet_leaf_6_wb_clk_i _02380_ _00683_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 _08013_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ clknet_leaf_53_wb_clk_i _02311_ _00614_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout492 _08025_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_6
X_13963_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08144__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10487__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ net1258 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
X_12914_ net365 _03612_ _03613_ net1054 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16682_ clknet_leaf_60_wb_clk_i _02242_ _00545_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_13894_ net1715 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[7\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__14217__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15633_ net1199 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
X_12845_ net2531 net215 net367 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ net2942 net254 net376 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ net1263 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ clknet_leaf_10_wb_clk_i _02863_ _01166_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14515_ net1317 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
X_11727_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\] _07023_ net675 vssd1 vssd1
+ vccd1 vccd1 _07868_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ net1181 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17234_ clknet_leaf_39_wb_clk_i _02794_ _01097_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14446_ net1384 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
X_11658_ net1674 net1157 net569 net1110 vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10609_ _05135_ _05099_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_107_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14377_ net1328 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
X_17165_ clknet_leaf_19_wb_clk_i _02725_ _01028_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10564__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08604__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ net1155 _04720_ _06844_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold907 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold918 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ net1404 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__inv_2
XANTENNA__12951__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13328_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _03745_ sky130_fd_sc_hd__and2_1
X_17096_ clknet_leaf_63_wb_clk_i _02656_ _00959_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold929 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ net1 net814 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nor2_2
X_16047_ net1368 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1607 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net3223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1618 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3234 sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ clknet_leaf_65_wb_clk_i _03547_ _01818_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3245 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17655__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09092__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16949_ clknet_leaf_9_wb_clk_i _02509_ _00812_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15391__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13904__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10031__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14208__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09421_ _05680_ _05682_ net575 _05654_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a31o_4
XFILLER_0_71_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09820__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09352_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] net618 _05586_
+ _05603_ _05607_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_87_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\]
+ net1046 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] net662 _05522_
+ _05529_ _05531_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14735__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout235_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08234_ net1683 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03513_ sky130_fd_sc_hd__mux2_1
XANTENNA__17035__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ net1711 net551 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1
+ vccd1 vccd1 _03530_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout402_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08452__B _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08096_ net1061 _04489_ _04492_ team_01_WB.instance_to_wrap.cpu.f0.i\[22\] _04518_
+ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09267__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17185__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1311_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09564__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout771_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout869_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] net867
+ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__and3_1
XANTENNA__10181__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12458__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13655__A0 _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10960_ _05487_ _06606_ _06608_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08908__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09874__A2 _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] net664 _05855_ _05859_
+ net670 vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a2111o_1
X_10891_ _05136_ _07154_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12630_ _08011_ _08017_ net488 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3_4
XFILLER_0_17_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ net2297 net295 net406 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08834__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] _07732_ _07753_ vssd1 vssd1 vccd1
+ vccd1 _07755_ sky130_fd_sc_hd__or3_1
X_14300_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\] _04444_ vssd1 vssd1 vccd1
+ vccd1 _04445_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09739__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15280_ net1257 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
X_12492_ net1875 net261 net413 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14231_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\] _04253_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a221o_1
X_11443_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] net1162 _04604_ _07683_ vssd1
+ vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16402__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08362__B _04624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12933__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\] _04246_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\]
+ _04311_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11374_ _07079_ _07629_ _07636_ _07637_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__a211o_1
X_13113_ net3084 _00017_ net357 _03726_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ _06578_ _06583_ _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14093_ net792 _04232_ _04243_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13044_ net1668 net834 net354 _03682_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a22o_1
X_17921_ clknet_leaf_101_wb_clk_i net2547 _01741_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09474__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16552__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17678__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _06516_ _06518_ _06519_ _06488_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__o31a_4
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1221 net1227 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17852_ clknet_leaf_77_wb_clk_i _03402_ _01672_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1232 net1235 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_4
XANTENNA__12104__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ net579 _06450_ _06416_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__o21a_1
XANTENNA__10413__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1243 net1245 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_4
Xfanout1254 net1261 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ clknet_leaf_132_wb_clk_i _02363_ _00666_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1265 net1267 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
Xfanout1276 net1301 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_2
Xfanout1287 net1289 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
X_17783_ clknet_leaf_113_wb_clk_i _03341_ _01604_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14995_ net1177 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
Xfanout1298 net1300 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__buf_4
XANTENNA__11943__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ clknet_leaf_139_wb_clk_i _02294_ _00597_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13946_ net1163 net1057 net3262 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[27\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11121__A1 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09640__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16665_ clknet_leaf_105_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[19\]
+ _00528_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13877_ net1159 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ _04142_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15616_ net1272 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12828_ _07842_ _08008_ net488 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16596_ clknet_leaf_57_wb_clk_i _02224_ _00459_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09617__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15547_ net1319 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
XANTENNA__08825__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12774__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ net2249 net296 net381 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15478_ net1303 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
X_17217_ clknet_leaf_129_wb_clk_i _02777_ _01080_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ net1233 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18197_ net1571 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
X_18076__1450 vssd1 vssd1 vccd1 vccd1 _18076__1450/HI net1450 sky130_fd_sc_hd__conb_1
XFILLER_0_13_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold704 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net2320
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17148_ clknet_leaf_12_wb_clk_i _02708_ _01011_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09087__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold726 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 _03506_ vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold748 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] net615 _06216_ _06222_
+ _06223_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__a2111o_1
Xhold759 team_01_WB.instance_to_wrap.cpu.f0.num\[5\] vssd1 vssd1 vccd1 vccd1 net2375
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ clknet_leaf_12_wb_clk_i _02639_ _00942_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10026__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08921_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] net887 vssd1
+ vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__and3_1
XANTENNA__13618__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08852_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] net842 vssd1
+ vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__and3_1
XANTENNA__12014__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1404 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11360__B2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1426 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _03440_ vssd1 vssd1 vccd1 vccd1 net3053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08783_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] net664 net638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\]
+ _05046_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a221o_1
Xhold1448 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1459 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13101__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13949__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] net896
+ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09335_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\] net851
+ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__and3_1
XANTENNA__12684__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14465__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09266_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\] net868 vssd1
+ vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__and3_1
XANTENNA__09559__A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14184__B _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08217_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_65_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09197_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] net851 vssd1
+ vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12915__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ net2349 net552 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1
+ vccd1 vccd1 _03547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10926__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1634_A team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15296__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08079_ net1366 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10110_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\] net610 _06351_ _06357_
+ _06366_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09294__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11090_ _06110_ net337 _07353_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__o21ba_1
XANTENNA__13528__B _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13876__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\] _04777_ _06286_
+ _06288_ _06300_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13340__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11351__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\] vssd1 vssd1 vccd1 vccd1
+ net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _02058_ vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold42 _02081_ vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _01976_ vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12859__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] vssd1 vssd1 vccd1 vccd1
+ net1680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold75 team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\] vssd1 vssd1 vccd1 vccd1
+ net1691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11763__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13800_ net2133 net782 _04099_ _04101_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__o22a_1
Xhold86 _01957_ vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\] vssd1 vssd1 vccd1 vccd1
+ net1713 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ net2420 net317 net467 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
X_14780_ net1385 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
XANTENNA__11103__A1 _06869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ _04048_ _04045_ net783 net1806 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ _05043_ _05099_ _05166_ _05241_ net516 net502 vssd1 vssd1 vccd1 vccd1 _07207_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09460__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16450_ clknet_leaf_107_wb_clk_i net2813 _00313_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13662_ _03775_ _03791_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ net535 _07137_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15401_ net1214 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ net2495 net280 net397 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12594__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16381_ clknet_leaf_29_wb_clk_i _02015_ _00249_ vssd1 vssd1 vccd1 vccd1 team_01_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
X_13593_ _07926_ _03932_ net189 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17350__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18120_ net1494 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
X_12544_ net3106 net219 net404 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15332_ net1224 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08373__A _04624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16918__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18051_ net1613 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15263_ net1293 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12475_ net2702 net227 net411 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10408__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17002_ clknet_leaf_43_wb_clk_i _02562_ _00865_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12906__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ _07686_ net1866 _07685_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__mux2_1
X_14214_ _04153_ net487 _04368_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__or4_1
XANTENNA_6 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15194_ net1265 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17836__D net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14145_ net789 _04231_ _04237_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a32o_1
XANTENNA__11938__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net543 _07473_ _07080_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\] net919 vssd1
+ vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14076_ net791 _04236_ _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__and3_4
X_11288_ _06030_ _07198_ _06916_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09635__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ _04847_ net571 _03666_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17904_ clknet_leaf_101_wb_clk_i net3166 _01724_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_10239_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] net878 vssd1
+ vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10145__A2 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_2
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
XFILLER_0_20_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1062 team_01_WB.instance_to_wrap.cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1 net1062
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ clknet_leaf_87_wb_clk_i _00006_ _01656_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11893__A2 _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1073 net1076 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_1
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_2
XANTENNA__13454__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13095__A1 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17766_ clknet_leaf_97_wb_clk_i net2221 _01587_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14978_ net1290 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
XANTENNA__09838__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16717_ clknet_leaf_20_wb_clk_i _02277_ _00580_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09370__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13929_ net1165 net1059 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[10\] sky130_fd_sc_hd__and3b_1
X_17697_ clknet_leaf_71_wb_clk_i _03257_ _01536_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16448__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16648_ clknet_leaf_88_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[2\]
+ _00511_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13901__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ clknet_leaf_123_wb_clk_i _02207_ _00442_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\] net908 vssd1
+ vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] net877
+ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__and3_1
XANTENNA__17843__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12009__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold501 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold512 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\] vssd1 vssd1 vccd1 vccd1
+ net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11848__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08577__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13570__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11581__A1 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17993__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\] vssd1 vssd1 vccd1 vccd1
+ net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\] vssd1 vssd1 vccd1 vccd1
+ net2205 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] net865 vssd1
+ vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13322__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] net668 vssd1 vssd1
+ vccd1 vccd1 _05168_ sky130_fd_sc_hd__or2_1
XANTENNA__10053__A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10136__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] net862 vssd1
+ vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1107_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09842__A _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1212 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] net762 _05097_ _05098_
+ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11884__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12679__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1234 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1 vccd1
+ net2850 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1245 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\] vssd1 vssd1 vccd1 vccd1
+ net2861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout567_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13086__A1 _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\] net700 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\]
+ _05021_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a221o_1
Xhold1278 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 net137 vssd1 vssd1 vccd1 vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08458__A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08697_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] net944 vssd1
+ vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout734_A _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17373__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__A0 _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09289__A _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ _06844_ _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09249_ _05502_ _05506_ _05510_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__or4_4
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ net2465 net261 net437 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__mux2_1
XANTENNA__13010__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11758__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ net520 net509 _06966_ _07472_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__o31a_1
XANTENNA__08568__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12191_ net2447 net317 net443 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__mux2_1
XANTENNA__10375__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _07404_ _07405_ net529 vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
X_15950_ net1395 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__inv_2
X_11073_ _07273_ _07333_ _07336_ _07085_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__o31a_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
X_10024_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] net899 vssd1
+ vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__and3_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ net1186 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12589__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ net1357 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__inv_2
XANTENNA__08740__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17620_ clknet_leaf_6_wb_clk_i _03180_ _01483_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14832_ net1346 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
XANTENNA__13077__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17716__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14274__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_101_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17551_ clknet_leaf_18_wb_clk_i _03111_ _01414_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09190__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14763_ net1246 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XANTENNA__11627__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ net2507 net230 net469 vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__mux2_1
XANTENNA_output117_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16502_ clknet_leaf_80_wb_clk_i net2776 _00365_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_13714_ net564 _04023_ _04033_ _04034_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17482_ clknet_leaf_41_wb_clk_i _03042_ _01345_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ net542 _07171_ _07080_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14694_ net1378 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XANTENNA__16740__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17866__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16433_ clknet_leaf_99_wb_clk_i _02061_ _00296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\]
+ sky130_fd_sc_hd__dfstp_1
X_13645_ net187 _07964_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
X_10857_ _06868_ _06950_ _06987_ _07083_ _07120_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__o41a_4
XANTENNA__10850__A3 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09199__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16364_ clknet_leaf_65_wb_clk_i net1850 _00232_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_140_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08307__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10788_ _06752_ _06697_ net499 vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__mux2_1
X_13576_ _03918_ _03917_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] net966
+ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09453__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10704__C_N _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ net1477 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ net1186 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
X_12527_ net2966 net307 net410 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16295_ clknet_leaf_113_wb_clk_i _01929_ _00163_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ net1600 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
X_15246_ net1228 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
XANTENNA__09205__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net2506 net301 net417 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08559__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ _07671_ _07672_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15177_ net1212 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
X_12389_ net2095 net304 net424 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
XANTENNA__10366__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14128_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\] _04239_ _04246_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\]
+ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a22o_1
XANTENNA__09365__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14059_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] _04221_ net566 vssd1
+ vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_24_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10118__A2 _06381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10304__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12499__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16270__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] net650 net627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17396__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17818_ clknet_leaf_67_wb_clk_i _03375_ _01639_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08731__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14265__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _04812_ _04813_ _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__or3_1
XANTENNA__08709__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17749_ clknet_leaf_116_wb_clk_i _03307_ _01570_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08482_ net1114 net1111 net1108 net1106 vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__and4b_4
XFILLER_0_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10747__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13240__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09103_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] net746 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13791__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09034_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] net705 _05283_
+ _05285_ _05287_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1057_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold320 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold331 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold342 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08460__B net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\] vssd1 vssd1 vccd1 vccd1
+ net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 _03746_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout684_A _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold397 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net815 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08970__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09936_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] net952 vssd1
+ vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__and3_1
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10109__A2 _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 _03727_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout844 _04772_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_8
Xfanout866 _04752_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
XANTENNA_fanout851_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] net736 _06116_ _06119_
+ _06121_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__a2111o_1
Xfanout877 _04746_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_4
Xfanout888 _04742_ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_2
Xhold1020 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\] vssd1 vssd1 vccd1 vccd1
+ net2636 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 net902 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
Xhold1031 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\] vssd1 vssd1 vccd1 vccd1
+ net2647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 team_01_WB.instance_to_wrap.a1.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2658
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1053 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 net2669
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12202__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\] net729 net695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09798_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] net734 _06045_ _06052_
+ _06053_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a2111o_1
Xhold1064 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16763__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] vssd1 vssd1 vccd1 vccd1
+ net2713 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17889__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _04988_ _05011_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11760_ net774 _07862_ _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08916__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _06697_ _06643_ net498 vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11691_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__nand2_1
XFILLER_0_95_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13430_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _06415_ vssd1 vssd1 vccd1
+ vccd1 _03783_ sky130_fd_sc_hd__and2_1
X_10642_ _05651_ _05686_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08789__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13361_ net24 net802 _03747_ net2252 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a22o_1
X_10573_ _06723_ _06777_ _06835_ _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__o31ai_1
XANTENNA__12872__S net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15100_ net1277 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ net3098 net221 net428 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__mux2_1
XANTENNA__09747__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13292_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] _04508_ team_01_WB.instance_to_wrap.a1.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__and3b_1
X_16080_ net1376 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__inv_2
XANTENNA__08651__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15031_ net1244 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
X_12243_ net2148 net228 net435 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13534__A2 _07640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11545__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11545__B2 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12174_ net2326 net233 net445 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11125_ _05378_ _05448_ _05515_ _05583_ net503 net518 vssd1 vssd1 vccd1 vccd1 _07389_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08961__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16982_ clknet_leaf_33_wb_clk_i _02542_ _00845_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12901__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10124__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15933_ net1342 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__inv_2
X_11056_ _07269_ _07277_ net524 vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10505__C1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10007_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\] net719 net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\]
+ _06256_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__a221o_1
XANTENNA__13208__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15864_ net1256 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__inv_2
XANTENNA__12112__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14247__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17603_ clknet_leaf_119_wb_clk_i _03163_ _01466_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14815_ net1384 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15795_ net1188 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__inv_2
XANTENNA__11951__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13732__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17534_ clknet_leaf_12_wb_clk_i _03094_ _01397_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14746_ net1293 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13470__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11958_ net2065 net242 net473 vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13451__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10909_ net520 _07172_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__and2_1
X_17465_ clknet_leaf_14_wb_clk_i _03025_ _01328_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14677_ net1369 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XANTENNA__10823__A3 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11889_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] net778 _07999_ _08000_
+ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_39_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16416_ clknet_leaf_103_wb_clk_i _02044_ _00279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_89_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ net770 _03961_ net969 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a21oi_1
X_17396_ clknet_leaf_4_wb_clk_i _02956_ _01259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16347_ clknet_leaf_64_wb_clk_i net1718 _00215_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13773__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12782__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13559_ _03845_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09657__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16278_ clknet_leaf_71_wb_clk_i _01915_ _00146_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09729__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18017_ net1594 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15229_ net1282 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09095__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15394__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10034__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _05981_ _05982_ _05983_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__or4_1
XANTENNA__16786__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09823__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13118__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _05912_ _05913_ _05914_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__or4_1
XANTENNA__12022__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14238__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08603_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\] net699 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a22o_1
X_09583_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] net733 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout265_A _07967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08534_ net549 _04796_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08465_ net996 net910 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__and2_4
XANTENNA_fanout432_A _08023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1174_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ net974 net935 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and2_1
XANTENNA__09417__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11224__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12692__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12972__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout899_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11527__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17561__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 _03446_ vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold161 team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] vssd1 vssd1 vccd1 vccd1
+ net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 net78 vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _03497_ vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1 vccd1
+ net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 _04764_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_8
Xfanout641 _04757_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_4
X_09919_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] net736 net698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__a22o_1
Xfanout652 _04745_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_8
Xfanout663 _04734_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_8
XANTENNA__09733__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_4
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_8
X_12930_ net1026 _07223_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__nand2_1
Xfanout696 _04688_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10241__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14229__B1 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12861_ team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] team_01_WB.instance_to_wrap.cpu.RU0.state\[2\]
+ net1059 net1165 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__o31a_1
XFILLER_0_115_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14600_ net1408 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11812_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] net676 net776 vssd1 vssd1
+ vccd1 vccd1 _07938_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15580_ net1234 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12792_ net2161 net296 net378 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XANTENNA__16509__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08646__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13452__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14531_ net1318 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
X_11743_ _07864_ _07880_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__nor2_1
XANTENNA__08864__D1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17250_ clknet_leaf_143_wb_clk_i _02810_ _01113_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14462_ net1392 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11674_ net2517 net1159 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16201_ clknet_leaf_95_wb_clk_i _01868_ _00069_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13413_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] _06773_ vssd1 vssd1
+ vccd1 vccd1 _03766_ sky130_fd_sc_hd__nand2_1
X_10625_ _06178_ _06179_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__nor2_1
X_17181_ clknet_leaf_127_wb_clk_i _02741_ _01044_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14393_ net1380 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11766__A1 _07324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16132_ net1321 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17904__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13344_ net12 net801 net596 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1
+ vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a22o_1
X_10556_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] net658 net624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\]
+ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__a221o_1
XANTENNA__08381__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__C _04644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16063_ net1368 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__inv_2
X_13275_ net1769 net810 net597 team_01_WB.instance_to_wrap.a1.ADR_I\[16\] vssd1 vssd1
+ vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
XANTENNA__10416__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__o21a_1
XANTENNA__12107__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ net1275 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
X_12226_ net2207 net298 net442 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__mux2_1
XANTENNA__12191__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11946__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13727__A _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ net2881 net304 net448 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11108_ _06041_ _06899_ _07371_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__o21a_1
X_12088_ net2074 net268 net458 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
X_16965_ clknet_leaf_134_wb_clk_i _02525_ _00828_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09643__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15916_ net1381 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__inv_2
X_11039_ _06856_ _06867_ _07302_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__and3_1
X_16896_ clknet_leaf_2_wb_clk_i _02456_ _00759_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09940__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15847_ net1195 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__inv_2
XANTENNA__12777__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13462__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15778_ net1290 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17434__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09151__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17517_ clknet_leaf_53_wb_clk_i _03077_ _01380_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14729_ net1320 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] net1798 net1047 vssd1 vssd1
+ vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
X_17448_ clknet_leaf_45_wb_clk_i _03008_ _01311_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08870__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ _04575_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__nor2_1
XANTENNA__15389__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17379_ clknet_leaf_120_wb_clk_i _02939_ _01242_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17584__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10029__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12954__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09818__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12017__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09178__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14171__A2 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08925__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] net951
+ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__and3_1
XANTENNA__15852__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10061__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09850__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09350__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\] net927
+ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12687__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1291_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A _04751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1389_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] net915 vssd1
+ vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08466__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09102__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\] net650 net632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\]
+ _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout814_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09497_ _05758_ _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16801__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08448_ _04703_ _04704_ _04709_ _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08379_ net1124 net953 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__and2_2
X_10410_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] net956
+ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09297__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11390_ _07082_ _07585_ _07611_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__and3b_1
XFILLER_0_34_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _06602_ _06603_ _06038_ _06044_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__a211o_2
XFILLER_0_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _05276_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__o21a_1
XANTENNA__09169__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10272_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] net895 vssd1
+ vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__and3_1
XANTENNA__14162__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__S net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ net2712 net227 net463 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17307__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1403 net1404 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1414 net1415 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 _08015_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout471 _08010_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ clknet_leaf_56_wb_clk_i _02310_ _00613_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15762__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 _07847_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_8
X_13962_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__and4bb_1
Xfanout493 _08025_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10487__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15701_ net1177 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_79_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12913_ net1031 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] vssd1 vssd1 vccd1
+ vccd1 _03613_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16681_ clknet_leaf_60_wb_clk_i _02241_ _00544_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13893_ net2320 net797 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_57_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15632_ net1262 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
X_12844_ net2054 net280 net368 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08807__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15563_ net1205 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ net2809 _07925_ net375 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ clknet_leaf_32_wb_clk_i _02862_ _01165_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ net1345 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
X_11726_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] _07866_ vssd1 vssd1
+ vccd1 vccd1 _07867_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15494_ net1287 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17233_ clknet_leaf_22_wb_clk_i _02793_ _01096_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14445_ net1385 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11657_ net3119 net1158 net569 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1
+ vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11739__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11530__A team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13221__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17164_ clknet_leaf_46_wb_clk_i _02724_ _01027_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10608_ _05015_ _05069_ _05138_ _05206_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__and4b_1
XFILLER_0_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ net1328 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XANTENNA__09638__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11588_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] _07807_ net840 vssd1 vssd1
+ vccd1 vccd1 _07808_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_107_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16115_ net1400 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__inv_2
XANTENNA__08542__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13327_ net1652 net808 net803 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold908 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\] vssd1 vssd1 vccd1 vccd1
+ net2524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold919 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\] net725 _06781_
+ _06786_ _06790_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_29_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17095_ clknet_leaf_130_wb_clk_i _02655_ _00958_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14153__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16046_ net1373 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__inv_2
X_13258_ team_01_WB.instance_to_wrap.a1.curr_state\[2\] team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13361__B1 _03747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12209_ net2707 net199 net439 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__mux2_1
X_13189_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
Xhold1608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3224 sky130_fd_sc_hd__dlygate4sd3_1
X_17997_ clknet_leaf_65_wb_clk_i _03546_ _01817_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13113__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16948_ clknet_leaf_4_wb_clk_i _02508_ _00811_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13904__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ clknet_leaf_54_wb_clk_i _02439_ _00742_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16824__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09420_ _05673_ _05674_ _05675_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__nor4_1
XANTENNA__12300__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\] net612 _05593_ _05597_
+ _05602_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11427__B1 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ net2647 net2508 net1041 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] net650 _05517_
+ _05521_ net670 vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16974__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ net1721 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout228_A _07911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08164_ net1777 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1
+ vccd1 vccd1 _03531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16204__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08095_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _04491_ _04493_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__o22a_1
XANTENNA__12970__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10056__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1137_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__A _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14144__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13352__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1304_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08997_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] net903
+ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11666__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09618_ _05878_ _05879_ _05880_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__or4_2
XANTENNA__12210__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _06607_ _06610_ _05138_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09549_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\] net644 _05793_ _05798_
+ _05802_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_136_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ net3074 net310 net406 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__mux2_1
XANTENNA__08834__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18169__1543 vssd1 vssd1 vccd1 vccd1 _18169__1543/HI net1543 sky130_fd_sc_hd__conb_1
XFILLER_0_52_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11511_ net483 _07753_ net319 vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ net2351 net300 net414 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\] _04268_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ _07696_ net1945 _07685_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_126_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09458__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12394__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13976__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15757__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14161_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\] _04233_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\]
+ _04310_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ _06955_ _07281_ _07336_ _07001_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ _06584_ _06585_ _06586_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__or4_1
X_13112_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\] _06559_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__mux2_1
XANTENNA_input60_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14135__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] _04252_ _04253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\]
+ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11496__S team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13343__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\] _03681_ net1029 vssd1
+ vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__mux2_1
X_10255_ _06508_ _06509_ _06510_ _06511_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ clknet_leaf_101_wb_clk_i net2874 _01740_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1203 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_2
Xfanout1211 net1236 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_2
X_17851_ clknet_leaf_80_wb_clk_i _03401_ _01671_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] net667 _06446_ _06449_
+ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__o22a_4
Xfanout1222 net1227 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09193__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18125__1499 vssd1 vssd1 vccd1 vccd1 _18125__1499/HI net1499 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
XFILLER_0_100_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1244 net1245 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
Xfanout1255 net1261 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_2
X_16802_ clknet_leaf_143_wb_clk_i _02362_ _00665_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08770__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17782_ clknet_leaf_113_wb_clk_i _03340_ _01603_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1266 net1267 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_4
Xfanout1277 net1285 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_4
XANTENNA__13646__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14994_ net1174 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XANTENNA__10132__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 net293 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_2
Xfanout1288 net1289 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_2
Xfanout1299 net1300 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09314__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16733_ clknet_leaf_126_wb_clk_i _02293_ _00596_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13945_ net1163 net1057 net3263 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[26\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__11657__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11121__A2 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13216__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12120__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ clknet_leaf_105_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[18\]
+ _00527_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13876_ net1165 net2521 net1055 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a21o_1
XANTENNA__16997__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15615_ net1294 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08537__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ net2637 net214 net374 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16595_ clknet_leaf_65_wb_clk_i _02223_ _00458_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15546_ net1305 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
X_12758_ net2609 net308 net381 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ _07849_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15477_ net1179 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12689_ net3064 net301 net389 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17216_ clknet_leaf_2_wb_clk_i _02776_ _01079_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14428_ net1234 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18196_ net1570 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
XFILLER_0_25_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09368__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17147_ clknet_leaf_32_wb_clk_i _02707_ _01010_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold705 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12790__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14359_ net1382 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09250__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10396__B1 _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold716 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10307__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold727 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09665__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ clknet_leaf_29_wb_clk_i _02638_ _00941_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold749 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16029_ net1355 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__inv_2
X_08920_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] net865
+ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__and3_1
XANTENNA__10604__A _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09553__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\] net882
+ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1405 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3043 sky130_fd_sc_hd__dlygate4sd3_1
X_08782_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] net652 net616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a22o_1
Xhold1438 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net3054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1449 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09305__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13126__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10320__B1 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09403_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\] net842
+ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout345_A _06870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\] net881
+ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\] net871
+ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout512_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1254_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__or4b_1
X_09196_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\] net863
+ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ net1697 net551 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1
+ vccd1 vccd1 _03548_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10387__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ net1 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__inv_2
XANTENNA__09792__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10139__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] net651 _06283_ _06292_
+ _06302_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold10 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[6\] vssd1 vssd1 vccd1 vccd1 net1626
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13247__D _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 team_01_WB.instance_to_wrap.a1.ADR_I\[4\] vssd1 vssd1 vccd1 vccd1 net1637
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\] vssd1 vssd1 vccd1 vccd1
+ net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\] vssd1 vssd1 vccd1 vccd1
+ net1659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold54 team_01_WB.instance_to_wrap.a1.ADR_I\[7\] vssd1 vssd1 vccd1 vccd1 net1670
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _03511_ vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold76 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\] vssd1 vssd1 vccd1 vccd1
+ net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net1703 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09741__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11991_ net2160 net304 net468 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
Xhold98 _03518_ vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11345__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ net786 _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ _05309_ _05378_ _05448_ _05515_ net503 net516 vssd1 vssd1 vccd1 vccd1 _07206_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10311__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08357__C net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13661_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] _03989_ net1067 vssd1
+ vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10873_ _07032_ _07036_ net530 vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15400_ net1207 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12612_ net2367 net251 net396 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16380_ clknet_leaf_112_wb_clk_i net1754 _00248_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13592_ _03925_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15331_ net1223 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12543_ net3135 net282 net403 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08373__B _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18050_ net1612 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
X_15262_ net1297 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12474_ net3132 net198 net411 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09188__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17001_ clknet_leaf_40_wb_clk_i _02561_ _00864_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17645__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ _04360_ _04361_ _04369_ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11425_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] net1162 vssd1 vssd1 vccd1
+ vccd1 _07686_ sky130_fd_sc_hd__and2_1
X_15193_ net1191 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XANTENNA_7 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10127__C _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\] _04247_ _04272_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\]
+ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__a221o_1
XANTENNA__14108__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11356_ _07618_ _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11590__A2 _07809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] net946 vssd1
+ vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12115__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14075_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__and2b_2
XFILLER_0_123_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17795__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ _06869_ _07536_ _07537_ _07550_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__a31o_2
XFILLER_0_120_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13026_ _03668_ _03669_ net355 net836 net1738 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a32o_1
X_17903_ clknet_leaf_107_wb_clk_i _03453_ _01723_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10238_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\] net886 vssd1
+ vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11954__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11342__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1041 net1046 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_4
X_10169_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] net883 vssd1
+ vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__and3_1
Xfanout1052 team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1 vccd1 net1052
+ sky130_fd_sc_hd__clkbuf_4
X_17834_ clknet_leaf_87_wb_clk_i _00016_ _01655_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout1063 team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1 vccd1 vccd1 net1063
+ sky130_fd_sc_hd__buf_2
XFILLER_0_94_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10550__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1074 net1076 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_2
Xfanout1085 net1088 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 net1105 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__buf_2
X_14977_ net1286 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
X_17765_ clknet_leaf_88_wb_clk_i _03323_ _01586_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13095__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16716_ clknet_leaf_44_wb_clk_i _02276_ _00579_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13928_ net1167 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[9\] sky130_fd_sc_hd__and3b_1
X_17696_ clknet_leaf_71_wb_clk_i _03256_ _01535_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16647_ clknet_leaf_86_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[1\]
+ _00510_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13859_ net2237 _04118_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[13\]
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12785__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17175__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16578_ clknet_leaf_141_wb_clk_i _02206_ _00441_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15529_ net1206 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] net892
+ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13555__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18179_ net1553 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
XFILLER_0_25_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold502 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10037__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold513 _02067_ vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09395__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold546 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09826__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13307__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold568 _02075_ vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12025__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\] net884 vssd1
+ vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08903_ net1113 net764 _04849_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__a21o_1
XANTENNA__11149__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] net865 vssd1
+ vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__and3_1
XANTENNA__10053__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18168__1542 vssd1 vssd1 vccd1 vccd1 _18168__1542/HI net1542 sky130_fd_sc_hd__conb_1
XANTENNA__13645__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] net710 net758 vssd1
+ vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__o21a_1
Xhold1213 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\] vssd1 vssd1 vccd1 vccd1
+ net2829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1002_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\] vssd1 vssd1 vccd1 vccd1
+ net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 _03399_ vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1246 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\] vssd1 vssd1 vccd1 vccd1
+ net2862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\] vssd1 vssd1 vccd1 vccd1
+ net2873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09561__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] net725 _05016_
+ _05022_ _05025_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13086__A2 _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_A _08015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1268 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
X_08696_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] net935 vssd1
+ vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10844__A1 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12695__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1371_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17668__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _05571_ _05575_ _05580_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__or3_4
XFILLER_0_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08905__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18124__1498 vssd1 vssd1 vccd1 vccd1 _18124__1498/HI net1498 sky130_fd_sc_hd__conb_1
X_09248_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\] net700 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\]
+ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09179_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\] net742 net726 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a22o_1
XANTENNA__16692__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11210_ _06991_ _07473_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__or2_1
X_12190_ net2335 net302 net444 vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09736__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08973__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ _07356_ _07359_ net513 vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__mux2_1
XANTENNA__10780__A0 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17048__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__09517__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ net532 net521 _07096_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__and3_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
X_10023_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\] net905 vssd1
+ vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__and3_1
X_14900_ net1258 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XANTENNA__11774__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08725__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15880_ net1357 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__inv_2
XANTENNA__08649__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ net1346 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13077__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08368__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17550_ clknet_leaf_53_wb_clk_i _03110_ _01413_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11088__A1 _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14762_ net1230 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
X_11974_ net2405 net236 net467 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__mux2_1
X_16501_ clknet_leaf_78_wb_clk_i net2543 _00364_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10410__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ team_01_WB.instance_to_wrap.cpu.f0.i\[28\] _04028_ _04029_ vssd1 vssd1 vccd1
+ vccd1 _04034_ sky130_fd_sc_hd__o21ba_1
X_17481_ clknet_leaf_42_wb_clk_i _03041_ _01344_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ _07187_ _07188_ net526 vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__mux2_1
X_14693_ net1375 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16432_ clknet_leaf_106_wb_clk_i _02060_ _00295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11803__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13644_ _03802_ _03970_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_141_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08384__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ net508 _06985_ _07117_ _07119_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08815__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16363_ clknet_leaf_68_wb_clk_i net1735 _00231_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13575_ net773 _07196_ net966 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__a21o_1
XANTENNA__09453__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ _04988_ _06807_ net499 vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__mux2_1
X_18102_ net1476 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__11014__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15314_ net1178 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
X_12526_ net2307 net313 net410 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
X_16294_ clknet_leaf_112_wb_clk_i _01928_ _00162_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11949__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18033_ net1599 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
X_15245_ net1214 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ net2396 net243 net417 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16106__A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11408_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _06486_ _06487_ vssd1
+ vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__or3_1
XANTENNA__13939__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15176_ net1181 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
X_12388_ net2623 net262 net424 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14127_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] _04287_ vssd1 vssd1 vccd1
+ vccd1 _04288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11339_ _05067_ _07290_ net346 vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__o21a_1
XANTENNA__10154__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ _04221_ net565 _04220_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and3b_1
X_13009_ net2246 net304 net362 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XANTENNA__13465__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17817_ clknet_leaf_67_wb_clk_i _03374_ _01638_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15680__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\] net742 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a22o_1
X_17748_ clknet_leaf_115_wb_clk_i _03306_ _01569_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17810__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08481_ net1070 net882 vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and2_4
X_17679_ clknet_leaf_74_wb_clk_i _03239_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11713__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13776__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09102_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] net728 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11251__B2 _07185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] net692 _05288_
+ _05292_ net712 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout308_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11003__B2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold321 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\] vssd1 vssd1 vccd1 vccd1
+ net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08460__C net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold354 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10064__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold365 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 team_01_WB.instance_to_wrap.cpu.c0.count\[8\] vssd1 vssd1 vccd1 vccd1 net1992
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1217_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09853__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold398 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _03745_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_4
Xfanout812 net815 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_2
XFILLER_0_106_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09935_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] net696 _06197_ _06198_
+ net713 vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__a2111o_1
Xfanout823 net833 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_2
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout677_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12503__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
Xfanout856 _04756_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
X_09866_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] net730 _06111_ _06123_
+ _06124_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a2111o_1
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
Xfanout878 _04746_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_4
Xhold1010 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\] vssd1 vssd1 vccd1 vccd1
+ net2626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net976 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] net961 vssd1
+ vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__and3_1
Xhold1032 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09291__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1043 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] net690 _06047_ _06049_
+ _06050_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__a2111o_1
Xhold1065 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08748_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__inv_2
Xhold1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10230__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17490__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] net658 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__inv_2
XANTENNA__10293__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ net2477 _07837_ net34 vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _05718_ _05753_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10045__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ net27 net802 _03747_ net1790 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XANTENNA__08643__C1 _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ _06665_ _06720_ _06667_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13519__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ net2317 net282 net427 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
X_13291_ net1853 net812 net597 team_01_WB.instance_to_wrap.a1.ADR_I\[0\] vssd1 vssd1
+ vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15030_ net1260 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
X_12242_ net2680 net199 net435 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__mux2_1
XANTENNA__09466__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16438__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ net3037 net234 net443 vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10405__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ _07386_ _07387_ net529 vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__mux2_1
X_16981_ clknet_leaf_8_wb_clk_i _02541_ _00844_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15932_ net1342 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__inv_2
X_11055_ _07314_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__nand2_1
XANTENNA__10702__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08379__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\] _04667_ net690 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\]
+ _06250_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a221o_1
X_15863_ net1238 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17833__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17602_ clknet_leaf_144_wb_clk_i _03162_ _01465_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14814_ net1357 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15794_ net1175 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__inv_2
X_14745_ net1277 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
X_17533_ clknet_leaf_14_wb_clk_i _03093_ _01396_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ net2245 net314 net472 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13224__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17983__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17464_ clknet_leaf_25_wb_clk_i _03024_ _01327_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ net514 _06966_ _07168_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14676_ net1373 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
X_11888_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\] net677 net778 vssd1 vssd1
+ vccd1 vccd1 _08000_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16415_ clknet_leaf_76_wb_clk_i _02043_ _00278_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13758__B1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ net770 _07551_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__or2_1
X_17395_ clknet_leaf_50_wb_clk_i _02955_ _01258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10839_ _06989_ _07102_ _07100_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18167__1541 vssd1 vssd1 vccd1 vccd1 _18167__1541/HI net1541 sky130_fd_sc_hd__conb_1
X_16346_ clknet_leaf_63_wb_clk_i net1817 _00214_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09938__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13558_ _03853_ _03902_ _03848_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21a_1
XANTENNA__17213__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12509_ net2551 net224 net408 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
X_16277_ clknet_leaf_71_wb_clk_i _01914_ _00145_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13489_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _05010_ vssd1 vssd1
+ vccd1 vccd1 _03842_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15228_ net1277 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
X_18016_ net107 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15159_ net1246 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10744__A0 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09673__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13907__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] net697 _05968_
+ _05976_ _05978_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11708__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12303__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18123__1497 vssd1 vssd1 vccd1 vccd1 _18123__1497/HI net1497 sky130_fd_sc_hd__conb_1
X_09651_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] net698 _05900_
+ _05901_ _05907_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09901__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08602_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\] net921 vssd1
+ vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__and3_1
X_09582_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] net727 net718 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09114__B1 _05376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ net549 _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ net1106 net1108 net1111 net1114 vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__nor4_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08455__C net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10059__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08395_ net1147 net1149 net1151 net1153 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout425_A _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1167_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09848__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08752__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12972__B2 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14174__B1 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ _05241_ _05277_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 net128 vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15585__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold151 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\] vssd1 vssd1 vccd1 vccd1
+ net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _01995_ vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold184 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16730__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 team_01_WB.instance_to_wrap.cpu.f0.write_data\[25\] vssd1 vssd1 vccd1 vccd1
+ net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout961_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 _04770_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_6
Xfanout631 _04763_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_6
X_09918_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\] net744 _04676_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__a22o_1
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12213__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 _04743_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_6
XANTENNA__11824__A1_N net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 _04732_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08156__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout675 net680 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_2
Xfanout686 _04695_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_6
XFILLER_0_77_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09849_ net1146 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] net949 vssd1
+ vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__and3_1
Xfanout697 _04687_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_6
XANTENNA__11160__B1 _06869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08561__D1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12860_ net2379 net212 net369 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09105__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ net676 _07520_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ net2847 net309 net378 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14530_ net1318 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XANTENNA__10266__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _07863_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13979__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14461_ net1336 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
X_11673_ net1820 net1159 net569 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1
+ vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ clknet_leaf_94_wb_clk_i _01867_ _00068_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_13412_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10624_ _06319_ _06887_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nand2_1
X_17180_ clknet_leaf_14_wb_clk_i _02740_ _01043_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14392_ net1380 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16131_ net1395 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13343_ net14 net798 net593 net2683 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17386__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] net910 vssd1
+ vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08631__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14165__B1 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16062_ net1374 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__inv_2
X_13274_ net1967 net812 net597 team_01_WB.instance_to_wrap.a1.ADR_I\[17\] vssd1 vssd1
+ vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
XANTENNA__09196__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ _06741_ _06742_ _06746_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__or4_2
X_15013_ net1225 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12225_ net2696 net242 net441 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__mux2_1
XANTENNA__10135__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net2675 net262 net448 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11107_ _06041_ _06899_ net324 vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12123__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16964_ clknet_leaf_13_wb_clk_i _02524_ _00827_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12087_ net2287 net272 net455 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_1
XANTENNA__08147__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15915_ net1387 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__inv_2
X_11038_ _06876_ _07159_ _05069_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16895_ clknet_leaf_1_wb_clk_i _02455_ _00758_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11962__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18011__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15846_ net1274 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__inv_2
XANTENNA__08837__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ net1313 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__inv_2
X_12989_ net2957 net208 net361 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ clknet_leaf_44_wb_clk_i _03076_ _01379_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14728_ net1331 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12793__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14659_ net1347 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
X_17447_ clknet_leaf_126_wb_clk_i _03007_ _01310_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10009__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ _04552_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\] team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__or3b_2
X_17378_ clknet_leaf_144_wb_clk_i _02938_ _01241_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16329_ clknet_leaf_63_wb_clk_i net1873 _00197_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08622__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14156__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17879__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09583__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12033__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__A _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] net961
+ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\] net938
+ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__and3_1
XANTENNA__10496__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12890__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17259__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\] net950 vssd1
+ vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout542_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08466__B net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1284_A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\] net639 net635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09496_ _05718_ _05753_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__xor2_4
XFILLER_0_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08447_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] net747 net713 _04698_
+ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout807_A _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08861__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire306 _07599_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08378_ net1149 net1153 net1151 net1148 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_74_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08913__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12208__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08613__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ _06602_ _06603_ _06044_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10271_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\] net884 vssd1
+ vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09574__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ net2753 net200 net463 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
XANTENNA__13370__B2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09744__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1404 net1413 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1415 net38 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 _08019_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 _08015_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 _08010_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _04154_
+ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18166__1540 vssd1 vssd1 vccd1 vccd1 _18166__1540/HI net1540 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 _07702_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09877__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout494 _07844_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12912_ net1027 _07287_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__nand2_1
X_15700_ net1240 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XANTENNA__13563__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16680_ clknet_leaf_61_wb_clk_i _02240_ _00543_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10487__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12881__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13892_ net2808 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[5\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_115_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15631_ net1249 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
X_12843_ net1845 net251 net370 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16626__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15562_ net1197 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12774_ net2032 net284 net377 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ net1345 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ clknet_leaf_8_wb_clk_i _02861_ _01164_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11725_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _07865_ vssd1 vssd1
+ vccd1 vccd1 _07866_ sky130_fd_sc_hd__nand2_1
X_15493_ net1229 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11811__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ net1395 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XANTENNA__09488__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17232_ clknet_leaf_25_wb_clk_i _02792_ _01095_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ net3018 net1157 net567 net1098 vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16776__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08392__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11739__A2 _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17163_ clknet_leaf_51_wb_clk_i _02723_ _01026_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12936__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18122__1496 vssd1 vssd1 vccd1 vccd1 _18122__1496/HI net1496 sky130_fd_sc_hd__conb_1
X_10607_ _04799_ _06842_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__or2_1
X_14375_ net1382 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08604__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _06847_ _04720_ vssd1 vssd1
+ vccd1 vccd1 _07807_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_10_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14138__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16114_ net1402 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13326_ net107 net814 net599 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ _06791_ _06799_ _06800_ _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__or4_1
X_17094_ clknet_leaf_141_wb_clk_i _02654_ _00957_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold909 _02126_ vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16045_ net1347 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__inv_2
X_13257_ team_01_WB.instance_to_wrap.a1.curr_state\[2\] team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10469_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\] net938
+ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12208_ net3144 net287 net439 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__mux2_1
XANTENNA__13361__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ net2699 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\] net820 vssd1 vssd1
+ vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11258__A _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ net2959 net204 net449 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
XANTENNA__10162__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17996_ clknet_leaf_56_wb_clk_i _03545_ _01816_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3225 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09951__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16947_ clknet_leaf_50_wb_clk_i _02507_ _00810_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12788__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10478__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12872__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16878_ clknet_leaf_55_wb_clk_i _02438_ _00741_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15829_ net1176 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__inv_2
XANTENNA__11705__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09350_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] net648 _05585_ _05592_
+ net671 vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17551__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08301_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\] net1765 net1044 vssd1 vssd1
+ vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ _05541_ _05542_ _05543_ _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11721__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ net1038 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09829__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ net1691 net551 net348 net1064 vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12028__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14129__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ _04477_ team_01_WB.instance_to_wrap.cpu.f0.num\[8\] team_01_WB.instance_to_wrap.cpu.f0.num\[10\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09556__B1 _05789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09564__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11363__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] net897 vssd1
+ vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__and3_1
XANTENNA__13104__A1 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14301__B1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12698__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout757_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16649__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11666__B2 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09617_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\] net609 _05860_ _05861_
+ _05876_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08908__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout924_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09548_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\] net634 _05791_ _05800_
+ _05805_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] net618 _05724_
+ _05733_ _05737_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08834__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11510_ _07718_ _07739_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12490_ net2834 net242 net413 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XANTENNA__09739__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ _04601_ _07683_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__a22o_1
XANTENNA__12918__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14160_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\] _04244_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\]
+ _04309_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a221o_1
XANTENNA__09795__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ _07054_ _07635_ _07632_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08940__A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13111_ net1746 net837 net357 _03725_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10323_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] net694 _06561_ _06570_
+ _06573_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14091_ net791 _04232_ _04236_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16179__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13042_ _06772_ net571 net359 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__o21a_1
XANTENNA_input53_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] net611 _06517_ net673
+ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__a211o_1
XANTENNA__17424__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09474__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_4
X_17850_ clknet_leaf_78_wb_clk_i _03400_ _01670_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10185_ _06440_ _06441_ _06447_ _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1223 net1227 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__buf_4
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_4
XANTENNA__10413__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16801_ clknet_leaf_138_wb_clk_i _02361_ _00664_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1245 net1268 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_2
Xfanout1256 net1261 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
X_17781_ clknet_leaf_116_wb_clk_i _03339_ _01602_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1267 net1268 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__clkbuf_4
Xfanout1278 net1285 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
XANTENNA__14389__A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
X_14993_ net1200 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
Xfanout291 net293 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1289 net1301 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17574__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ clknet_leaf_20_wb_clk_i _02292_ _00595_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13944_ net1163 net1057 net3261 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[25\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__12401__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13875_ net1166 net1060 net1625 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a21o_1
X_16663_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[17\]
+ _00526_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11017__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ net2523 net291 net372 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
X_15614_ net1292 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09078__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16594_ clknet_leaf_68_wb_clk_i _02222_ _00457_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ net3239 net312 net381 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15545_ net1190 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XANTENNA__08825__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11541__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13232__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _07848_ vssd1 vssd1 vccd1
+ vccd1 _07849_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ net1241 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12688_ net2203 net245 net390 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14427_ net1234 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
X_17215_ clknet_leaf_1_wb_clk_i _02775_ _01078_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11639_ net1835 net1797 net840 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__mux2_1
X_18195_ net1569 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13582__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14358_ net3207 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__clkbuf_1
X_17146_ clknet_leaf_33_wb_clk_i _02706_ _01009_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ net1730 net809 net804 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\] vssd1
+ vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
Xhold728 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17077_ clknet_leaf_9_wb_clk_i _02637_ _00940_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold739 team_01_WB.instance_to_wrap.cpu.f0.num\[31\] vssd1 vssd1 vccd1 vccd1 net2355
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14289_ _04194_ _04438_ _04201_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__o21a_1
X_16028_ net1410 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__inv_2
XANTENNA_wire558_A _05751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08210__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08850_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\] net860
+ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17917__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09681__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1406 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net3022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1417 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3033 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] net635 net626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\]
+ _05044_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a221o_1
X_17979_ clknet_leaf_70_wb_clk_i _03528_ _01799_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1428 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1439 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3055 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11716__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16941__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] net847 vssd1
+ vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\] net867
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13270__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11451__A team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout338_A _06983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] net882 vssd1
+ vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09195_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\] net868
+ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1247_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08146_ net1685 net551 net348 net1061 vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a22o_1
XANTENNA__09856__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16321__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09241__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08077_ team_01_WB.instance_to_wrap.a1.READ_I vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1414_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09294__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08201__A0 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1522_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17597__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10233__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\] vssd1 vssd1 vccd1 vccd1
+ net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 _01987_ vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[3\] vssd1 vssd1 vccd1 vccd1 net1649
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\] vssd1 vssd1 vccd1 vccd1
+ net1660 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _04627_ net764 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__or2_1
Xhold55 _01990_ vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 net89 vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] vssd1 vssd1 vccd1 vccd1
+ net1693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12221__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 net110 vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net3137 net263 net470 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
X_18121__1495 vssd1 vssd1 vccd1 vccd1 _18121__1495/HI net1495 sky130_fd_sc_hd__conb_1
Xhold99 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net1715
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10847__C1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _05756_ _07203_ _05622_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__a21o_1
X_13660_ net769 _03987_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _07076_ _07135_ _07079_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ net2778 net256 net397 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13261__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ _03834_ _03924_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13800__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15330_ net1311 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XANTENNA__11967__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12542_ net2767 net223 net405 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09480__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15261_ net1281 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XANTENNA__15768__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12891__S net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ net3161 net286 net411 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17000_ clknet_leaf_62_wb_clk_i _02560_ _00863_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10408__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14212_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\] _04266_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ _04364_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__a221o_1
X_11424_ _04503_ _07683_ _07684_ _07681_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09766__A _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13564__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15192_ net1257 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
XANTENNA_8 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14143_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] _04258_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\]
+ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11355_ net521 _07019_ _07185_ _07576_ _06971_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__a32o_1
XANTENNA__08440__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10306_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] net959 vssd1
+ vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__and3_1
X_14074_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__and2_2
XFILLER_0_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11286_ _07200_ _07539_ _07540_ _07549_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11327__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ net837 team_01_WB.instance_to_wrap.cpu.RU0.next_write_i vssd1 vssd1 vccd1
+ vccd1 _03670_ sky130_fd_sc_hd__and2b_1
X_17902_ clknet_leaf_99_wb_clk_i _03452_ _01722_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] net846 vssd1
+ vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1031 net1036 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_2
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
X_17833_ clknet_leaf_87_wb_clk_i _00015_ _01654_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10168_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\] net909 vssd1
+ vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__and3_1
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
XANTENNA__16964__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 net1064
+ sky130_fd_sc_hd__buf_2
XANTENNA__11536__A team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_94_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_1
Xfanout1086 net1088 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_2
XANTENNA__15008__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17764_ clknet_leaf_88_wb_clk_i _03322_ _01585_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1097 net1098 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_2
X_10099_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] net888 vssd1
+ vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__and3_1
X_14976_ net1269 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_63_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16715_ clknet_leaf_51_wb_clk_i _02275_ _00578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13927_ net1165 net1059 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[8\] sky130_fd_sc_hd__and3b_1
X_17695_ clknet_leaf_84_wb_clk_i _03255_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11970__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16646_ clknet_leaf_88_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[0\]
+ _00509_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13858_ _04118_ _04137_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08845__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12809_ net2837 net254 net372 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16577_ clknet_leaf_129_wb_clk_i _02205_ _00440_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13789_ net1064 net1065 _07705_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1
+ vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15528_ net1197 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15678__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15459_ net1223 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
XANTENNA__13555__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09676__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18178_ net1552 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
X_18145__1519 vssd1 vssd1 vccd1 vccd1 _18145__1519/HI net1519 sky130_fd_sc_hd__conb_1
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold503 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ clknet_leaf_40_wb_clk_i _02689_ _00992_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16494__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold514 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\] vssd1 vssd1 vccd1 vccd1
+ net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12306__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__A _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold536 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\] vssd1 vssd1 vccd1 vccd1
+ net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\] net848 vssd1
+ vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__and3_1
Xhold558 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08902_ net560 _05165_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] net762
+ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\] net899 vssd1
+ vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and3_1
XANTENNA__10714__A_N _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ _05087_ _05089_ _05093_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or4_2
Xhold1203 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout190_A _07874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1225 _02046_ vssd1 vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1236 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12041__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] net950
+ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__and3_1
Xhold1258 _03470_ vssd1 vssd1 vccd1 vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
X_08695_ _04957_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout455_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__S net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1197_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08755__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout622_A _04768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1364_A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ _05576_ _05577_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__or4_1
XANTENNA__09998__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09247_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] net697 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__a22o_1
XANTENNA__08670__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16837__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10228__C net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09178_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] net733 _05439_ _05440_
+ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09214__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout991_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08921__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08129_ _04503_ _04555_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or2_4
XFILLER_0_82_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12216__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ _07357_ _07403_ net517 vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__mux2_1
XANTENNA__16987__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10780__A1 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _07273_ _07333_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__nor2_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
X_10022_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] net873 vssd1
+ vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16217__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1347 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
XANTENNA__14274__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14761_ net1216 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
X_11973_ net2430 net202 net469 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16500_ clknet_leaf_102_wb_clk_i net2529 _00363_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_13712_ net1061 _04022_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__or2_1
X_10924_ _06961_ _07006_ net510 vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__mux2_1
X_17480_ clknet_leaf_45_wb_clk_i _03040_ _01343_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14692_ net1400 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16431_ clknet_leaf_77_wb_clk_i _02059_ _00294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13234__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13643_ net968 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _03974_ _03975_
+ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
X_10855_ _07116_ _07118_ _07099_ _07103_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08384__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16362_ clknet_leaf_65_wb_clk_i net1914 _00230_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
X_13574_ net186 _07912_ _03916_ net767 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__o211a_1
XANTENNA__09199__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ _07046_ _07049_ net525 vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__mux2_1
XANTENNA__10599__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09453__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18101_ net1475 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_109_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15313_ net1246 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
X_12525_ net2045 net261 net410 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
X_16293_ clknet_leaf_98_wb_clk_i _01927_ _00161_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18032_ net1426 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XANTENNA__09496__A _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12456_ net2875 net314 net416 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
X_15244_ net1266 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XANTENNA__09205__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11407_ _06486_ _06487_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1
+ vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15175_ net1183 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12387_ net2681 net268 net426 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__mux2_1
XANTENNA__12126__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14126_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] net789 vssd1 vssd1 vccd1
+ vccd1 _04287_ sky130_fd_sc_hd__nand2_1
X_11338_ _05067_ net344 _07290_ _07601_ _05015_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__o311a_1
XFILLER_0_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10771__A1 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ _04218_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and3_1
X_11269_ _07107_ _07531_ _07532_ _07529_ _07530_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__o311a_1
X_13008_ net1909 net264 net362 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
XANTENNA__09662__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17142__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11266__A _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17816_ clknet_leaf_67_wb_clk_i _03373_ _01637_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14265__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17747_ clknet_leaf_106_wb_clk_i _03305_ _01568_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12796__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ net1201 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13481__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ net1106 net1108 net1111 net1114 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__and4bb_2
X_17678_ clknet_leaf_73_wb_clk_i _03238_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__17292__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09692__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16629_ clknet_leaf_104_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[15\]
+ _00492_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11713__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13776__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09444__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] _04680_ _05355_
+ _05357_ _05359_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09032_ _05290_ _05293_ _05294_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120__1494 vssd1 vssd1 vccd1 vccd1 _18120__1494/HI net1494 sky130_fd_sc_hd__conb_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold300 _01994_ vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12036__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold311 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout203_A _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10211__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold333 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 net1971
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold388 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 _03745_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_106_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold399 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\] net931 vssd1
+ vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__and3_1
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1112_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout824 net833 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__buf_2
XFILLER_0_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_2
Xfanout857 _04756_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_2
X_09865_ _06126_ _06127_ _06128_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__or3_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 _04750_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
Xhold1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 _04746_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_4
Xhold1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\] net916
+ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__and3_1
Xhold1044 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\] vssd1 vssd1 vccd1 vccd1
+ net2660 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] net719 _04696_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1055 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 net2693
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _05009_ _05010_ net580 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__mux2_1
Xhold1088 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net2704
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1099 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\] vssd1 vssd1 vccd1 vccd1
+ net2715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout837_A _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08678_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\] net652 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\]
+ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a221o_1
XANTENNA__08485__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08916__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17785__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10640_ _06900_ _06902_ _06903_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _06776_ _06830_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__and2b_1
XANTENNA__11242__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ net2865 net224 net429 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10450__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ net86 net812 net597 net1801 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XANTENNA__17015__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09747__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08651__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12241_ net2532 net288 net435 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14950__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ net2852 net203 net445 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11785__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17165__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11123_ net548 _05718_ _05923_ _05993_ net504 net518 vssd1 vssd1 vccd1 vccd1 _07387_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16980_ clknet_leaf_9_wb_clk_i _02540_ _00843_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ net1342 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__inv_2
X_11054_ net321 _07317_ _07311_ _07002_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08379__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] _04651_ _06266_
+ _06267_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a2111o_1
X_15862_ net1304 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14247__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17601_ clknet_leaf_137_wb_clk_i _03161_ _01464_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14813_ net1352 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
X_15793_ net1192 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
X_18144__1518 vssd1 vssd1 vccd1 vccd1 _18144__1518/HI net1518 sky130_fd_sc_hd__conb_1
XFILLER_0_19_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17532_ clknet_leaf_14_wb_clk_i _03092_ _01395_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14744_ net1277 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
X_11956_ net2319 net302 net474 vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ net537 _07069_ _07170_ _07166_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a31o_1
X_17463_ clknet_leaf_11_wb_clk_i _03023_ _01326_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11887_ net678 _07456_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14675_ net1361 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16414_ clknet_leaf_83_wb_clk_i _02042_ _00277_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10838_ _07101_ net338 _06593_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13626_ _07950_ _03960_ net188 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__mux2_1
X_17394_ clknet_leaf_31_wb_clk_i _02954_ _01257_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16345_ clknet_leaf_63_wb_clk_i net1757 _00213_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08634__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13557_ _03841_ _03850_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__and2_1
X_10769_ _07029_ _07032_ net528 vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__mux2_1
XANTENNA__16117__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15021__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12508_ net2548 net226 net407 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
X_16276_ clknet_leaf_66_wb_clk_i _01913_ _00144_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13488_ _03836_ _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18015_ net107 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15227_ net1299 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
X_12439_ net2915 net230 net415 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17508__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08937__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09954__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ net1259 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10744__A1 _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\] _04266_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\]
+ _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__a221o_1
X_15089_ net1189 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17658__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09650_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\] net694 _05893_
+ _05899_ _05905_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14238__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\] net941
+ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and3_1
XANTENNA__12249__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] net746 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\]
+ _05828_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a221o_1
XANTENNA__09114__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _04727_ _04795_ net583 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08463_ _04723_ _04726_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1
+ vccd1 vccd1 _04727_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17038__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08394_ net970 net940 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__and2_1
XANTENNA__09417__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08625__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12972__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10432__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ _05241_ _05277_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__or2_1
XANTENNA__17188__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15866__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1327_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 net1746
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _01979_ vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold152 _02123_ vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold163 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold174 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net1790
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_01_WB.instance_to_wrap.a1.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 net1801
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold196 team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\] vssd1 vssd1 vccd1 vccd1
+ net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _04776_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_8
Xfanout621 _04770_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout632 _04763_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_8
X_09917_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] net747 net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout643 _04755_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_8
Xfanout654 _04743_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13685__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 _04732_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_4
XANTENNA__10499__B1 _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net680 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_4
X_09848_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] net927 vssd1
+ vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and3_1
Xfanout687 _04693_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_8
Xfanout698 _04687_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10241__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14229__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ _05788_ _05822_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _07856_ _07935_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__or2_1
X_12790_ net2206 net313 net378 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09656__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11741_ net2996 net208 net481 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__mux2_1
XANTENNA__08646__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14460_ net1392 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
X_11672_ net1644 net1159 net568 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1
+ vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10623_ _06385_ _06456_ _06883_ _06886_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13411_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] _06773_ vssd1 vssd1
+ vccd1 vccd1 _03764_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12412__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14391_ net1380 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XANTENNA__16405__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16130_ net1394 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13342_ net15 net801 net596 net1665 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a22o_1
XANTENNA__10423__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\] net642 net638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\]
+ _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13273_ net1837 net812 net598 team_01_WB.instance_to_wrap.a1.ADR_I\[18\] vssd1 vssd1
+ vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
XANTENNA__14165__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15776__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ net1355 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10485_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\] net736 net713 _06747_
+ _06748_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_126_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15012_ net1271 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
X_12224_ net2560 net314 net439 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux2_1
XANTENNA__10416__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17800__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__B _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net2296 net268 net449 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__mux2_1
XANTENNA__12404__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _06602_ _06603_ _06041_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__a21o_1
X_16963_ clknet_leaf_131_wb_clk_i _02523_ _00826_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12086_ net2139 net247 net455 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15914_ net1387 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__inv_2
X_11037_ _07002_ _07294_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16894_ clknet_leaf_3_wb_clk_i _02454_ _00757_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17950__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15845_ net1232 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__inv_2
XANTENNA__09940__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11544__A team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15776_ net1273 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ net3215 net190 net360 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17515_ clknet_leaf_60_wb_clk_i _03075_ _01378_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09014__A _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14727_ net1314 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11939_ net2928 net234 net471 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__mux2_1
X_17446_ clknet_leaf_141_wb_clk_i _03006_ _01309_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14658_ net1409 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08853__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13609_ _03813_ _03820_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__and2_1
X_17377_ clknet_leaf_137_wb_clk_i _02937_ _01240_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14589_ net1376 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17330__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16328_ clknet_leaf_64_wb_clk_i net1705 _00196_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12954__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16259_ clknet_leaf_69_wb_clk_i net2585 _00127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17480__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11719__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10342__B _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] net917
+ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10061__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09633_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] net958
+ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09850__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout368_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__B2 _03596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__A team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09564_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] net957 vssd1
+ vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09099__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14092__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\] net661 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09495_ _05718_ _05754_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout535_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1277_A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09859__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\] net723 net706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08763__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ net976 net957 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__and2_4
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire318 _07367_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16578__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09297__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10236__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18143__1517 vssd1 vssd1 vccd1 vccd1 _18143__1517/HI net1517 sky130_fd_sc_hd__conb_1
XFILLER_0_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09594__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] net651 _06531_ _06532_
+ _06533_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11905__A0 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12224__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10184__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17973__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1405 net1412 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__buf_4
XFILLER_0_100_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 _08021_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 _08018_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_6
Xfanout462 _08015_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ _04148_ _04150_ _04151_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 _08010_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout484 _04556_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 _07844_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_1
XANTENNA__17203__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ net2467 net607 net589 _03611_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12881__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13891_ net1846 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[4\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12881__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15630_ net1231 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12842_ net2831 net257 net368 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14083__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15561_ net1221 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12773_ net1879 net224 net377 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17353__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ clknet_leaf_7_wb_clk_i _02860_ _01163_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14512_ net1361 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _07864_ vssd1 vssd1
+ vccd1 vccd1 _07865_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15492_ net1269 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ clknet_leaf_54_wb_clk_i _02791_ _01094_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14443_ net1390 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
X_11655_ net2779 net1157 net567 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1
+ vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11811__B _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08392__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17162_ clknet_leaf_48_wb_clk_i _02722_ _01025_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10606_ _06866_ _06868_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__or2_2
X_14374_ net1328 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
X_11586_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _06847_ _04720_ vssd1 vssd1
+ vccd1 vccd1 _07806_ sky130_fd_sc_hd__o21a_4
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09801__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ net1365 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13325_ net1 _03741_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nand2_1
X_10537_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\] net738 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17093_ clknet_leaf_129_wb_clk_i _02653_ _00956_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16044_ net1410 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__inv_2
X_13256_ team_01_WB.EN_VAL_REG net72 _03739_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
X_10468_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\] net945 vssd1
+ vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11539__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ net2572 net230 net441 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13187_ net2890 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\] net824 vssd1 vssd1
+ vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
X_10399_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net763 net590 vssd1 vssd1
+ vccd1 vccd1 _06663_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12138_ net2725 net239 net447 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__mux2_1
XANTENNA__11258__B _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17995_ clknet_leaf_61_wb_clk_i _03544_ _01815_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11973__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13113__A2 _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16946_ clknet_leaf_23_wb_clk_i _02506_ _00809_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12069_ net3083 net192 net455 vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09868__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09670__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16877_ clknet_leaf_21_wb_clk_i _02437_ _00740_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12872__A1 _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10883__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15828_ net1242 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11588__B1_N net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15759_ net1246 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
XANTENNA__14585__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08300_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\] net2061 net1039 vssd1 vssd1
+ vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09679__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\] net624 _05518_ _05523_
+ _05535_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__mux2_1
X_17429_ clknet_leaf_25_wb_clk_i _02989_ _01292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11721__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12309__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08162_ net1687 net551 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1
+ vccd1 vccd1 _03533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08093_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\] team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16870__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10056__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13352__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10353__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17226__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] net881
+ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout485_A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13664__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11115__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_A _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16250__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17376__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09616_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] net622 _05857_ _05874_
+ _05875_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11418__A2 _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] _04741_ _05796_
+ _05797_ _05804_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13812__B1 _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout917_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09589__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08493__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\] net664 net616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08429_ net1118 net913 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12219__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _07695_ net1939 _07685_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13040__A1 _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09244__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11371_ net525 _07315_ _07633_ _07634_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13110_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\] _06520_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__mux2_1
X_10322_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\] net717 net706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14090_ net790 net787 _04236_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__and3_4
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ net1847 net834 net355 _03680_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] net645 net613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__a22o_1
XANTENNA__13343__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__A1 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input46_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\] net617 _06420_ _06430_
+ _06436_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
Xfanout1213 net1218 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1224 net1227 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
X_16800_ clknet_leaf_142_wb_clk_i _02360_ _00663_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08770__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1249 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_4
X_17780_ clknet_leaf_116_wb_clk_i _03338_ _01601_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_135_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14992_ net1256 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
Xfanout1257 net1261 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_4
Xfanout1268 net1302 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_2
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout1279 net1285 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__buf_4
Xfanout281 _07939_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
X_16731_ clknet_leaf_39_wb_clk_i _02291_ _00594_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13943_ net1163 net1057 net2582 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[24\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08387__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08522__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10865__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16662_ clknet_leaf_104_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[16\]
+ _00525_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13874_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\] _04567_ team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en
+ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a21o_1
X_15613_ net1283 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XANTENNA__17869__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ net3040 net295 net374 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16593_ clknet_leaf_65_wb_clk_i _02221_ _00456_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13803__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15544_ net1255 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
X_12756_ net2587 net261 net381 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 _07848_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12129__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ net1188 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ net2511 net316 net387 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17214_ clknet_leaf_4_wb_clk_i _02774_ _01077_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14426_ net1279 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11638_ net1692 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] net840 vssd1 vssd1
+ vccd1 vccd1 _03323_ sky130_fd_sc_hd__mux2_1
X_18194_ net1568 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
XFILLER_0_25_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09235__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17145_ clknet_leaf_17_wb_clk_i _02705_ _01008_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14357_ net1781 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13582__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11569_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] net1161 vssd1 vssd1 vccd1 vccd1
+ _07794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10396__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire682 _04717_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_1
Xhold707 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ net115 net811 net806 net1622 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold718 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\] vssd1 vssd1 vccd1 vccd1
+ net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17076_ clknet_leaf_6_wb_clk_i _02636_ _00939_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09665__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14288_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\] _04193_ vssd1 vssd1 vccd1
+ vccd1 _04438_ sky130_fd_sc_hd__nor2_1
X_16027_ net1402 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13239_ _03723_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] net831 vssd1 vssd1
+ vccd1 vccd1 _02019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09962__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12799__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08780_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] net642 net610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a22o_1
Xhold1407 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\] vssd1 vssd1 vccd1 vccd1
+ net3023 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13098__A1 _06106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17978_ clknet_leaf_78_wb_clk_i _03527_ _01798_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1418 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3045 sky130_fd_sc_hd__dlygate4sd3_1
X_16929_ clknet_leaf_138_wb_clk_i _02489_ _00792_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10320__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\] net891 vssd1
+ vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18142__1516 vssd1 vssd1 vccd1 vccd1 _18142__1516/HI net1516 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09332_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\] net856 vssd1
+ vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__and3_1
XANTENNA__13270__A1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10084__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__B team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09202__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09263_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] net856
+ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout233_A _07897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12039__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08214_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09194_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] net891
+ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ net3180 net552 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1
+ vccd1 vccd1 _03550_ sky130_fd_sc_hd__a22o_1
XANTENNA__13659__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout400_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10387__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ team_01_WB.instance_to_wrap.a1.WRITE_I vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__inv_2
XANTENNA__08252__S net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15874__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16616__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1407_A net1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08201__A1 _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 net1628
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold23 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net1639
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__A1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] vssd1 vssd1 vccd1 vccd1
+ net1650 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net765 _04719_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1
+ vccd1 vccd1 _05242_ sky130_fd_sc_hd__o21a_1
Xhold45 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] vssd1 vssd1 vccd1 vccd1
+ net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\] vssd1 vssd1 vccd1 vccd1
+ net1683 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16766__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold78 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 net1694
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11626__B _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 _01962_ vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ _05756_ _07203_ _05622_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10311__A2 _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10871_ net537 _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ net2403 net220 net397 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ _03930_ _03929_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] net966
+ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ net2734 net226 net403 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ net1277 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ net2337 net231 net413 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08951__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14211_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\] _04260_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\]
+ _04365_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__a221o_1
X_11423_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04504_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\]
+ _04567_ _00019_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15191_ net1246 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11575__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10378__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__B2 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14142_ _04299_ _04300_ _04301_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11354_ _06955_ _07553_ _07617_ _05279_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] net922 vssd1
+ vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14073_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] _04227_ _04234_ vssd1 vssd1
+ vccd1 vccd1 _04235_ sky130_fd_sc_hd__a21o_1
X_11285_ net321 _07546_ _07548_ _07545_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__a211o_1
XANTENNA__17541__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10236_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] net868 vssd1
+ vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and3_1
X_13024_ _04510_ _03577_ _03580_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_write_i
+ sky130_fd_sc_hd__nor3b_1
XANTENNA__09782__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17901_ clknet_leaf_104_wb_clk_i _03451_ _01721_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_63_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 net1012 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_2
X_17832_ clknet_leaf_87_wb_clk_i _00005_ _01653_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10167_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] net869 vssd1
+ vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__and3_1
XANTENNA__12412__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1032 net1034 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__buf_2
Xfanout1043 net1046 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_1
XANTENNA__08398__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1065 team_01_WB.instance_to_wrap.cpu.f0.i\[7\] vssd1 vssd1 vccd1 vccd1 net1065
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10550__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11536__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17763_ clknet_leaf_88_wb_clk_i net2011 _01584_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1076 net1105 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12827__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_1
X_14975_ net1293 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
X_10098_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\] net906 vssd1
+ vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1098 net1105 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_4
X_16714_ clknet_leaf_49_wb_clk_i _02274_ _00577_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13926_ net1166 net1059 net1715 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[7\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17694_ clknet_leaf_84_wb_clk_i _03254_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16645_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[31\]
+ _00508_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13857_ net2424 _04117_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15024__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ net2984 net221 net372 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__mux2_1
X_16576_ clknet_leaf_129_wb_clk_i _02204_ _00439_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13788_ _07706_ _07780_ net484 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09022__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15527_ net1182 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_32_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ net2188 net226 net379 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09957__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ net1266 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XANTENNA__14201__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17071__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13555__A2 _07324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ net1309 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
X_18177_ net1551 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_0_89_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16639__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ net1281 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10369__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17128_ clknet_leaf_61_wb_clk_i _02688_ _00991_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold504 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold515 _03469_ vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09395__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold537 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\] vssd1 vssd1 vccd1 vccd1
+ net2164 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\] net908 vssd1
+ vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17059_ clknet_leaf_133_wb_clk_i _02619_ _00922_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold559 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08901_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] net710 net758 vssd1
+ vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__o21ai_1
X_09881_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\] net848 vssd1
+ vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and3_1
XANTENNA__08195__A0 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08832_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\] net717 net711 _05094_
+ _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12322__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1204 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\] vssd1 vssd1 vccd1 vccd1
+ net2820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14268__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] net940 vssd1
+ vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__and3_1
Xhold1259 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08694_ _04935_ _04956_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10844__A3 _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11462__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A _08019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08247__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17414__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] net748 _05556_
+ _05564_ _05566_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_118_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12992__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_A _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09246_ _05494_ _05507_ _05508_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08670__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] net746 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11557__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17564__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08128_ _04503_ _04555_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout984_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08059_ team_01_WB.instance_to_wrap.cpu.f0.num\[27\] vssd1 vssd1 vccd1 vccd1 _04490_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_124_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08973__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11070_ _07333_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__inv_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
X_10021_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\] net869 vssd1
+ vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__and3_1
XANTENNA__08725__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14259__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14760_ net1266 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
X_11972_ net2230 net239 net469 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13711_ net3250 net785 _04032_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09150__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10923_ _06956_ _06962_ net509 vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14691_ net1363 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16430_ clknet_leaf_80_wb_clk_i net1647 _00293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_13642_ net772 _07568_ net968 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10854_ _06991_ _06996_ net546 vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__a21o_1
XANTENNA__17094__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ clknet_leaf_65_wb_clk_i net1789 _00229_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
X_13573_ net186 _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__nand2_1
X_10785_ _07047_ _07048_ net516 vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__mux2_1
X_18100_ net1474 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
X_15312_ net1247 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
X_12524_ net2004 net300 net410 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
X_16292_ clknet_leaf_111_wb_clk_i _01926_ _00160_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18031_ net1425 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_15243_ net1210 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12455_ net2854 net302 net415 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12407__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ _07663_ _07668_ _04627_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__a21o_1
X_15174_ net1277 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ net2437 net272 net423 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08964__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14125_ net2036 net584 _04286_ net1170 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o211a_1
X_11337_ _06877_ _07302_ net322 vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18141__1515 vssd1 vssd1 vccd1 vccd1 _18141__1515/HI net1515 sky130_fd_sc_hd__conb_1
XFILLER_0_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12931__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10154__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14056_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04218_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11268_ net532 _07292_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007_ net2476 net268 net362 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
XANTENNA__08716__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ _06472_ _06474_ _06479_ _06482_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__or4_4
XFILLER_0_98_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12142__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ _06596_ _07458_ _07462_ _06972_ _07461_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11181__C1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17815_ clknet_leaf_68_wb_clk_i _03372_ _01636_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11981__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17746_ clknet_leaf_105_wb_clk_i _03304_ _01567_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14958_ net1230 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08856__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17437__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09141__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13909_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\] net794 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[22\] sky130_fd_sc_hd__and2_1
X_17677_ clknet_leaf_75_wb_clk_i _03237_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14889_ net1221 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16628_ clknet_leaf_104_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[14\]
+ _00491_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13225__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09429__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15689__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16559_ clknet_leaf_50_wb_clk_i _02187_ _00422_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16461__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09100_ _05361_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__or3_1
XANTENNA__12984__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08591__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09031_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] net742 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\]
+ _05282_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18229_ net601 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12317__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold301 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] vssd1 vssd1 vccd1 vccd1
+ net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold312 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\] vssd1 vssd1 vccd1 vccd1
+ net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[2\] vssd1 vssd1 vccd1 vccd1
+ net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold334 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _01971_ vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10064__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold367 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\] net938 vssd1
+ vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and3_1
Xhold389 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_2
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09853__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
Xfanout825 net833 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11457__A team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13148__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12052__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\] net704 net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a22o_1
XANTENNA__10361__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout847 _04769_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
Xfanout858 _04756_ vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_4
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_4
XANTENNA__11172__C1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\] vssd1 vssd1 vccd1 vccd1
+ net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] net949
+ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and3_1
XANTENNA__09380__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09795_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] net717 net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__a22o_1
XANTENNA__12987__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1034 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout565_A _04202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net2683
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] net763 net590 vssd1 vssd1
+ vccd1 vccd1 _05010_ sky130_fd_sc_hd__a21o_1
Xhold1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout732_A _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\] net662 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a22o_1
XANTENNA__08485__B net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16804__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11778__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09597__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10570_ _06723_ _06833_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__nor2_1
XANTENNA__08643__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16954__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09229_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\] net961
+ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12227__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ net2848 net230 net436 vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux2_1
XANTENNA__14192__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12171_ net2838 net239 net445 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
X_11122_ _05788_ _05852_ _06071_ _06141_ net504 net517 vssd1 vssd1 vccd1 vccd1 _07386_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold890 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
X_15930_ net1342 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__inv_2
X_11053_ _07312_ _07316_ net533 vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10505__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] _04645_ _06254_
+ _06258_ _06261_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09371__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ net1179 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17600_ clknet_leaf_2_wb_clk_i _03160_ _01463_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14812_ net1357 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09659__B1 _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15792_ net1244 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__inv_2
X_17531_ clknet_leaf_37_wb_clk_i _03091_ _01394_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1590 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14743_ net1317 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
X_11955_ net2526 net262 net472 vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__mux2_1
XANTENNA_output115_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ clknet_leaf_31_wb_clk_i _03022_ _01325_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10906_ net520 _07169_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14674_ net1409 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
X_11886_ net2955 net310 net482 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16413_ clknet_leaf_75_wb_clk_i _02041_ _00276_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13625_ _03819_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__xnor2_1
X_17393_ clknet_leaf_21_wb_clk_i _02953_ _01256_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10837_ _06867_ net342 vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12926__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16344_ clknet_leaf_64_wb_clk_i net1695 _00212_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XANTENNA__15302__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13556_ net967 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _03900_ _03901_
+ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ _07030_ _07031_ net518 vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__mux2_1
XANTENNA__09938__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ net2242 net199 net407 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
X_16275_ clknet_leaf_67_wb_clk_i _01912_ _00143_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12137__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _05244_ _03837_ _03839_
+ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_23_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10699_ _06961_ _06962_ net516 vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__mux2_1
X_18014_ net107 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
X_15226_ net1260 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
X_12438_ net3184 net234 net415 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11976__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13757__A team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08937__A2 _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15157_ net1177 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
X_12369_ net2191 net208 net425 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14108_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\] _04268_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09673__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15088_ net1257 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14039_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] _04147_ vssd1 vssd1 vccd1 vccd1
+ _04210_ sky130_fd_sc_hd__and4_1
XANTENNA__14013__A_N team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08600_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\] net925 vssd1
+ vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__and3_1
XANTENNA__13492__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08570__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16827__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ _05840_ _05841_ _05842_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__or4_1
XANTENNA__12600__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09114__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] net668 _04788_ _04794_
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__o22a_2
X_17729_ clknet_leaf_96_wb_clk_i _03287_ _01550_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08462_ net764 _04724_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ net1147 net1149 net1152 net1154 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__and4_4
XFILLER_0_50_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10059__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12957__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15212__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09848__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10432__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16207__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12047__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10356__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout313_A _07994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1055_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09014_ _05241_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__nand2_1
XANTENNA__14174__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11886__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold120 team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\] vssd1 vssd1 vccd1 vccd1
+ net1736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__A2 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1 vccd1
+ net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net124 vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 net82 vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16357__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\] vssd1 vssd1 vccd1 vccd1
+ net1791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08260__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 _01984_ vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] vssd1 vssd1 vccd1 vccd1
+ net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _03742_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
XFILLER_0_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout611 _04776_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_4
X_09916_ _06178_ _06179_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__nand2_1
Xfanout622 _04768_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10091__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout633 _04762_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_8
XFILLER_0_121_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_6
XANTENNA__13685__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 _04741_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_6
Xfanout666 net669 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_6
XANTENNA__09880__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] net954 vssd1
+ vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__and3_1
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_2
Xfanout688 _04693_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12510__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09778_ _05824_ _05891_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ _04989_ _04990_ _04991_ _04992_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__or4_1
XANTENNA__11634__B _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11740_ net774 _07876_ _07878_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_95_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18140__1514 vssd1 vssd1 vccd1 vccd1 _18140__1514/HI net1514 sky130_fd_sc_hd__conb_1
XFILLER_0_7_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ net2334 net1159 net568 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1
+ vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ _03761_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or2_1
XANTENNA__15122__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ _06385_ _06414_ net524 net536 _06347_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14390_ net1329 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13341_ net16 net798 net593 net3080 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__o22a_1
X_10553_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] net664 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16060_ net1410 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__inv_2
X_13272_ net85 net812 net598 net1775 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
XANTENNA__14165__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10484_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[25\] _04667_ _06727_
+ _06731_ _06736_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15011_ net1223 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12223_ net2052 net303 net440 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__mux2_1
XANTENNA__17282__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ net2811 net272 net447 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11105_ _06041_ _06602_ _06603_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nand3_1
X_12085_ net2079 net276 net456 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__mux2_1
XANTENNA__13676__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16962_ clknet_leaf_142_wb_clk_i _02522_ _00825_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09344__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15913_ net1383 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__inv_2
X_11036_ _07042_ _07185_ _07298_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16893_ clknet_leaf_130_wb_clk_i _02453_ _00756_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08552__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15844_ net1270 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__inv_2
XANTENNA__12420__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11439__B1 _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08837__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15775_ net1297 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12987_ net2684 net196 net361 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ clknet_leaf_42_wb_clk_i _03074_ _01377_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14726_ net1320 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11938_ net3198 net204 net473 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17445_ clknet_leaf_134_wb_clk_i _03005_ _01308_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14657_ net1399 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
X_11869_ net2949 net300 net481 vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__mux2_1
XANTENNA__09949__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13608_ net966 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _03944_ _03945_
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
X_17376_ clknet_leaf_142_wb_clk_i _02936_ _01239_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14588_ net1407 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16327_ clknet_leaf_57_wb_clk_i _01961_ _00195_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
X_13539_ net771 _07585_ _03885_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16258_ clknet_leaf_69_wb_clk_i _01895_ _00126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09965__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14156__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15209_ net1212 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16189_ clknet_leaf_91_wb_clk_i _01856_ _00057_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09583__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11719__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08791__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17775__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] net922 vssd1
+ vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13934__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09632_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\] net954 vssd1
+ vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and3_1
XANTENNA__12330__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12890__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17005__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09563_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\] net944 vssd1
+ vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout263_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08514_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\] net649 net645 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__a22o_1
X_09494_ net548 _05686_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__xor2_2
X_08445_ _04705_ _04706_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout430_A _08024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11470__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A _06451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08376_ net1150 net1151 net1153 net1148 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__nor4b_1
XANTENNA__08255__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1378_A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14781__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10517__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09875__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13355__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09574__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1406 net1412 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 _08024_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 _08021_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout452 _08018_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11669__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _08010_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 _04556_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 _07810_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_2
X_12910_ net366 _03609_ _03610_ net1056 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a32o_1
XANTENNA__12240__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13890_ net1790 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[3\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12841_ net2282 net219 net368 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
XANTENNA__14083__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15560_ net1181 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
X_12772_ net2769 net228 net375 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XANTENNA__08954__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14511_ net1361 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\]
+ _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ net1221 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17230_ clknet_leaf_51_wb_clk_i _02790_ _01093_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ net1395 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11654_ net2470 net1157 net567 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1
+ vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a22o_1
XANTENNA__17648__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17161_ clknet_leaf_39_wb_clk_i _02721_ _01024_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ _06866_ _06868_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__nor2_2
X_14373_ net1327 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11585_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[31\] net573 vssd1 vssd1 vccd1
+ vccd1 _07805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16112_ net1377 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__inv_2
X_13324_ net1815 net813 net807 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[0\] vssd1
+ vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a22o_1
XANTENNA__14138__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09785__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\] net749 _06780_
+ _06783_ _06792_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a2111o_1
X_17092_ clknet_leaf_128_wb_clk_i _02652_ _00955_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13346__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16043_ net1401 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13255_ net73 net71 net74 _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12415__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] net920
+ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__and3_1
XANTENNA__16672__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17798__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ net2919 net234 net439 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13186_ net1902 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\] net818 vssd1 vssd1
+ vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
X_10398_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] net668 _06655_ _06661_
+ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__o22a_2
XFILLER_0_23_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08773__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ net2216 net208 net449 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_1
X_17994_ clknet_leaf_58_wb_clk_i _03543_ _01814_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10162__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17028__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16945_ clknet_leaf_21_wb_clk_i _02505_ _00808_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12068_ net2168 net194 net457 vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__mux2_1
XANTENNA__09951__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08525__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12150__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _07078_ _07271_ _07275_ _07282_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16876_ clknet_leaf_48_wb_clk_i _02436_ _00739_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09025__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15827_ net1186 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15758_ net1217 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ net1375 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15689_ net1213 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11290__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08230_ net1728 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\] net1040 vssd1 vssd1
+ vccd1 vccd1 _03517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17428_ clknet_leaf_4_wb_clk_i _02988_ _01291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10618__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08161_ net1744 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1
+ vccd1 vccd1 _03534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18211__1585 vssd1 vssd1 vccd1 vccd1 _18211__1585/HI net1585 sky130_fd_sc_hd__conb_1
XFILLER_0_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17359_ clknet_leaf_18_wb_clk_i _02919_ _01222_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11060__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] team_01_WB.instance_to_wrap.cpu.f0.num\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14129__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13337__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12325__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12560__A1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\] net872 vssd1
+ vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1018_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09308__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13664__B _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08516__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13156__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09615_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] net614 _05856_ _05866_
+ _05873_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12995__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1387_A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09546_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] net664 net657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11823__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout812_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\] net648 net612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\]
+ _05730_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08493__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\] net925
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12379__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13576__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08359_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\] _04621_ vssd1 vssd1 vccd1 vccd1
+ _04623_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09795__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ net515 _07052_ net520 vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10321_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] net724 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\]
+ _06569_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12235__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13040_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\] _03679_ net1028 vssd1
+ vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09547__A2 _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ _06512_ _06513_ _06514_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__A2 _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10183_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\] net645 _06432_ _06438_
+ net673 vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__a2111o_1
Xfanout1203 net1302 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_2
XANTENNA__08949__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1214 net1218 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
Xfanout1225 net1227 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_4
Xfanout1236 net1302 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_2
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1247 net1249 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_4
X_14991_ net1248 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
Xfanout260 _07989_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout1258 net1260 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
Xfanout271 _07957_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
Xfanout1269 net1272 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_4
Xfanout282 _07920_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
XANTENNA__17320__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16730_ clknet_leaf_36_wb_clk_i _02290_ _00593_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13942_ net1163 net1057 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[23\] sky130_fd_sc_hd__and3b_1
XFILLER_0_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout293 _08004_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09180__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ clknet_leaf_95_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[15\]
+ _00524_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13873_ team_01_WB.instance_to_wrap.cpu.DM0.dhit net1162 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en sky130_fd_sc_hd__and2_1
X_15612_ net1279 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
X_12824_ net3011 net307 net374 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
X_16592_ clknet_leaf_65_wb_clk_i _02220_ _00455_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_104_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15543_ net1247 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
XANTENNA__11822__B _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12755_ net2088 net299 net381 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ net495 _07845_ _07846_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__and3_1
X_15474_ net1178 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
X_12686_ net2265 net305 net388 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14425_ net1279 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
X_17213_ clknet_leaf_127_wb_clk_i _02773_ _01076_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_18193_ net1567 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
X_11637_ net2220 net840 _07808_ _07833_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12934__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10157__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17144_ clknet_leaf_27_wb_clk_i _02704_ _01007_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14356_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1
+ vccd1 _02242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11568_ net320 _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13319__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ net116 net812 net806 net1628 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold708 team_01_WB.instance_to_wrap.cpu.f0.num\[21\] vssd1 vssd1 vccd1 vccd1 net2324
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12790__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17075_ clknet_leaf_48_wb_clk_i _02635_ _00938_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold719 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\] net935
+ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__and3_1
X_14287_ _04201_ _04437_ net1367 vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12145__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ _07744_ _07746_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ net1394 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__inv_2
X_13238_ _03722_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] net829 vssd1 vssd1
+ vccd1 vccd1 _02020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11984__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16418__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__A2 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ net2979 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\] net828 vssd1 vssd1
+ vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XANTENNA__10553__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1408 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3024 sky130_fd_sc_hd__dlygate4sd3_1
X_17977_ clknet_leaf_70_wb_clk_i _03526_ _01797_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09681__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1419 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16928_ clknet_leaf_2_wb_clk_i _02488_ _00791_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16568__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16859_ clknet_leaf_37_wb_clk_i _02419_ _00722_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17813__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09400_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\] net856 vssd1
+ vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13931__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09331_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\] net843
+ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10629__A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13270__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11281__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\] net907
+ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09193_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] net845
+ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout226_A _07911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08144_ net1812 net552 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[30\] vssd1 vssd1
+ vccd1 vccd1 _03551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13659__B _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08760__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12055__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ net1161 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_114_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1135_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10792__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11894__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10544__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1302_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 _01968_ vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] net760 _05239_ _05240_
+ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a22o_4
Xhold24 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\] vssd1 vssd1 vccd1 vccd1 net1640
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\] vssd1 vssd1 vccd1 vccd1
+ net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] vssd1 vssd1 vccd1 vccd1
+ net1673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold68 _03513_ vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _01978_ vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17493__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ net526 _07059_ _07071_ _07132_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09529_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\] net903 vssd1
+ vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13261__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10075__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ net2573 net201 net403 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13549__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12471_ net3204 net234 net411 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XANTENNA__09217__A1 _05480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__A1_N _06992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14210_ _04356_ _04357_ _04366_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__or4_1
XFILLER_0_129_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11422_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\] _07682_ vssd1 vssd1 vccd1 vccd1
+ _07683_ sky130_fd_sc_hd__nor2_2
XFILLER_0_30_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15190_ net1258 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\] _04227_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\]
+ _04292_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11353_ _05277_ net334 net333 _07616_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08440__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10783__A0 _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10304_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] net914 vssd1
+ vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__and3_1
X_14072_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] _04229_ _04233_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\]
+ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11284_ net535 _07165_ _07547_ _07106_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11327__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08728__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\] net1029 vssd1 vssd1 vccd1
+ vccd1 _03669_ sky130_fd_sc_hd__or2_1
X_17900_ clknet_leaf_75_wb_clk_i net2946 _01720_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] net851 vssd1
+ vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1000 net1008 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1022 net1023 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_2
X_17831_ clknet_leaf_87_wb_clk_i _00014_ _01652_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10166_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] net848 vssd1
+ vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__and3_1
Xfanout1033 net1034 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16710__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17836__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 net1045 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1055 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1055 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
X_17762_ clknet_leaf_89_wb_clk_i _03320_ _01583_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_18210__1584 vssd1 vssd1 vccd1 vccd1 _18210__1584/HI net1584 sky130_fd_sc_hd__conb_1
Xfanout1077 net1080 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_2
X_14974_ net1316 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
X_10097_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\] net869 vssd1
+ vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__and3_1
Xfanout1088 net1096 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09689__D1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
X_16713_ clknet_leaf_40_wb_clk_i _02273_ _00576_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10838__A1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13925_ net1166 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[6\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[6\] sky130_fd_sc_hd__and3b_1
X_17693_ clknet_leaf_82_wb_clk_i _03253_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11833__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ _04117_ net2435 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[11\]
+ sky130_fd_sc_hd__nor2_1
X_16644_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[30\]
+ _00507_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09303__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08845__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ net2017 net284 net371 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13787_ _04091_ _04089_ net782 net1794 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_85_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16575_ clknet_leaf_119_wb_clk_i _02203_ _00438_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09456__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10999_ _07002_ _07252_ _07259_ _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__o211a_1
XANTENNA__11393__A_N _07324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15526_ net1275 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
X_12738_ net2630 net198 net379 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17216__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11979__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15457_ net1312 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
X_12669_ net3163 net235 net387 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14408_ net1309 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
XANTENNA__09759__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18176_ net1550 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_72_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08353__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15388_ net1270 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09676__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11566__A2 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14339_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1 vssd1 vccd1
+ vccd1 _02259_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16240__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17127_ clknet_leaf_119_wb_clk_i _02687_ _00990_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17366__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold505 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold516 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold538 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
X_17058_ clknet_leaf_143_wb_clk_i _02618_ _00921_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold549 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16009_ net1363 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__inv_2
X_08900_ _05152_ _05153_ _05158_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__nor4_1
XANTENNA__13495__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] net905 vssd1
+ vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12603__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08195__A1 _04592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08589__A _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16390__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\] net734 _05071_ _05076_
+ _05083_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_104_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1205 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] net944
+ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__and3_1
Xhold1238 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10829__A1 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ _04935_ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__and2_1
XANTENNA__09695__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13779__B1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09314_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\] net742 net702 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09998__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09245_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\] net701 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17709__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\] net751 net718 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08263__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ _04536_ _04550_ _04555_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] vssd1
+ vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10525__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09883__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] vssd1 vssd1 vccd1 vccd1 _04489_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_102_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17859__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__C1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12513__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\] net844 vssd1
+ vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16883__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11971_ net2277 net206 net469 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13710_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] _04024_ _04029_ _04031_ net785
+ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__a311o_1
XANTENNA__10296__A2 _06559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15125__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ net545 _06970_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14690_ net1406 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17239__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ net769 _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__nand2_1
X_10853_ _06971_ _07105_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16360_ clknet_leaf_66_wb_clk_i net1916 _00228_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11245__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ _03849_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10784_ _05378_ _05309_ net502 vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15311_ net1248 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12523_ net2241 net242 net409 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XANTENNA__16263__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16291_ clknet_leaf_98_wb_clk_i _01925_ _00159_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17389__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08661__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18030_ net1424 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
X_15242_ net1197 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
X_12454_ net2247 net263 net416 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ _07663_ _07668_ _04627_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__a21oi_2
X_15173_ net1226 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12385_ net2963 net248 net424 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
X_14124_ _04235_ _04245_ _04251_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or4_2
XFILLER_0_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11336_ net346 _07587_ net306 vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_104_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13519__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14055_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04218_ _04219_ vssd1
+ vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11828__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ net539 _07390_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__nor2_1
XANTENNA__12423__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10508__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ net1901 net272 net360 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
X_10218_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] net702 _06480_ _06481_
+ net712 vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a2111o_1
X_11198_ net523 _07019_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11181__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17814_ clknet_leaf_67_wb_clk_i _03371_ _01635_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10149_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10170__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17745_ clknet_leaf_105_wb_clk_i _03303_ _01566_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14957_ net1212 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ net1665 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[21\]
+ sky130_fd_sc_hd__and2_1
X_17676_ clknet_leaf_73_wb_clk_i _03236_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14888_ net1201 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16627_ clknet_leaf_104_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[13\]
+ _00490_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13839_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04113_ vssd1 vssd1 vccd1 vccd1
+ _04129_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10039__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__A0 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16558_ clknet_leaf_39_wb_clk_i _02186_ _00421_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08101__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08872__A _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15509_ net1174 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ clknet_leaf_85_wb_clk_i _02117_ _00352_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10995__B1 _07258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] net701 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18228_ net1589 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18159_ net1533 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold302 _03418_ vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold313 _03326_ vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold324 _03393_ vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold335 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold346 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold368 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] net750 _06193_ _06194_
+ _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_22_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold379 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12333__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10642__A _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout815 _03740_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_4
Xfanout826 net827 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09904__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] net690 _06113_ _06114_
+ _06125_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a2111o_1
Xfanout837 _00017_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_8
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_4
XANTENNA_fanout293_A _08004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _04756_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_2
X_08814_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\] net936
+ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__and3_1
Xhold1002 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] vssd1 vssd1 vccd1 vccd1
+ net2618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1024 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\] vssd1 vssd1 vccd1 vccd1
+ net2640 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] net754 net698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\]
+ _06051_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a221o_1
Xhold1035 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1046 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] net666 _04998_ _05008_
+ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__o22a_4
Xhold1057 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A _08015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\] vssd1 vssd1 vccd1 vccd1
+ net2695 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13164__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10278__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08676_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\] net643 net625 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\]
+ _04937_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10089__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08891__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17531__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12975__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11778__A2 _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12975__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08643__A2 _04902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14177__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09228_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] net921
+ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10450__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09159_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\] net951 vssd1
+ vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12170_ net2276 net206 net445 vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11121_ _06971_ _07042_ _07384_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12243__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold880 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08159__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11052_ _07279_ _07315_ net522 vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] net733 net714 _06257_
+ _06260_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_102_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15860_ net1241 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__inv_2
XANTENNA__08957__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__B1 _06995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17061__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ net1357 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XANTENNA__10698__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15791_ net1201 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__inv_2
Xhold1580 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3196 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16629__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17530_ clknet_leaf_36_wb_clk_i _03090_ _01393_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14742_ net1331 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
Xhold1591 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3207 sky130_fd_sc_hd__dlygate4sd3_1
X_11954_ net1947 net266 net473 vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10905_ _07071_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__nand2_1
X_14673_ net1400 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
X_17461_ clknet_leaf_8_wb_clk_i _03021_ _01324_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11885_ _04622_ _07995_ _07996_ _07997_ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16412_ clknet_leaf_103_wb_clk_i _02040_ _00275_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13624_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05720_ _03946_ vssd1
+ vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10836_ net505 _06592_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__and2_1
XANTENNA__09788__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17392_ clknet_leaf_23_wb_clk_i _02952_ _01255_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16779__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12926__B _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16343_ clknet_leaf_63_wb_clk_i net1848 _00211_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
X_13555_ net767 _07324_ net1066 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__o21a_1
X_10767_ _05788_ _05993_ net504 vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__mux2_1
XANTENNA__12418__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08634__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ net3162 net286 net407 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__mux2_1
X_16274_ clknet_leaf_66_wb_clk_i _01911_ _00142_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10441__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13486_ _03831_ _03835_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _05309_ _05241_ net502 vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__mux2_1
X_18013_ net107 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
X_15225_ net1237 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
X_12437_ net3199 net202 net417 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10729__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13391__B2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15156_ net1241 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ net2256 net192 net423 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09954__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ net787 _04232_ _04236_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__and3_4
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11319_ _06668_ _07569_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10462__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15087_ net1201 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XANTENNA__12153__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12299_ _07842_ net494 _08008_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__and3_4
XANTENNA__16159__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ _04147_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1
+ _04209_ sky130_fd_sc_hd__a31o_1
XANTENNA__09028__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11992__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15989_ net1381 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17554__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _04790_ _04791_ _04792_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__or4_1
X_17728_ clknet_leaf_96_wb_clk_i _03286_ _01549_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08461_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] _04628_ _04635_ vssd1 vssd1
+ vccd1 vccd1 _04725_ sky130_fd_sc_hd__and3_1
X_17659_ clknet_leaf_36_wb_clk_i _03219_ _01522_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10722__A2_N net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08392_ net973 net943 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__and2_4
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12957__B2 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12328__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08625__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14159__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10432__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _05244_ _05276_ net583 vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__mux2_2
XFILLER_0_108_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1048_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 _01964_ vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13382__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold121 team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\] vssd1 vssd1 vccd1 vccd1
+ net1737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold132 team_01_WB.instance_to_wrap.cpu.c0.count\[0\] vssd1 vssd1 vccd1 vccd1 net1748
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold143 _01975_ vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _01999_ vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11468__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12063__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold176 _03482_ vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1215_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 net603 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_2
Xhold187 team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] vssd1 vssd1 vccd1 vccd1
+ net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _04775_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_6
X_09915_ _06141_ _06175_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__xor2_2
Xfanout623 _04768_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_4
XANTENNA__12998__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout634 _04762_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
Xfanout645 _04753_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_8
XANTENNA__13685__A2 _07456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_6
X_18089__1463 vssd1 vssd1 vccd1 vccd1 _18089__1463/HI net1463 sky130_fd_sc_hd__conb_1
Xfanout667 net668 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_8
X_09846_ _06071_ _06108_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__nand2_1
XANTENNA__10499__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net680 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_2
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_6
X_09777_ _05890_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout842_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08728_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] net635 net626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09510__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08659_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\] net753 net744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08864__A2 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13622__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11670_ net1635 net1159 net568 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1
+ vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__B2 _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ _06879_ _06884_ _06385_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__o21a_1
XANTENNA__09401__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12238__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11142__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13340_ net17 net798 net593 net2232 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10423__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ _06809_ _06811_ _06813_ _06815_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13271_ net1827 net812 net597 team_01_WB.instance_to_wrap.a1.ADR_I\[20\] vssd1 vssd1
+ vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10483_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\] net744 net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_129_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15010_ net1311 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
X_12222_ net2795 net264 net440 vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input69_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17427__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ net2015 net248 net447 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11104_ _07347_ _07348_ net318 vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16961_ clknet_leaf_136_wb_clk_i _02521_ _00824_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12084_ net1993 net217 net455 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13676__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15912_ net1387 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__inv_2
X_11035_ _06955_ _07033_ _07050_ _06971_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__a22o_1
XANTENNA__16451__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ clknet_leaf_11_wb_clk_i _02452_ _00755_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15843_ net1219 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ net1315 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12986_ net494 _07846_ _08011_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ clknet_leaf_41_wb_clk_i _03073_ _01376_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ net1322 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11937_ net2092 net239 net473 vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__mux2_1
XANTENNA__13532__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17444_ clknet_leaf_128_wb_clk_i _03004_ _01307_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14656_ net1402 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
X_11868_ net779 _07981_ _07982_ _07983_ vssd1 vssd1 vccd1 vccd1 _07984_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12939__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08853__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ net549 _04796_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__and2b_1
X_13607_ net768 _03943_ net967 vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12148__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17375_ clknet_leaf_1_wb_clk_i _02935_ _01238_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14587_ net1407 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
XANTENNA__08607__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\] net680 net775 vssd1 vssd1
+ vccd1 vccd1 _07927_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16326_ clknet_leaf_63_wb_clk_i net1762 _00194_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ net185 _03886_ net771 vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a21o_1
XANTENNA__09280__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11987__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16257_ clknet_leaf_69_wb_clk_i _01894_ _00125_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13469_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _05653_ _05720_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15208_ net1181 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16188_ clknet_leaf_91_wb_clk_i _01855_ _00056_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15139_ net1220 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\] net915 vssd1
+ vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12611__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__B1 _03584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13934__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09631_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\] net945 vssd1
+ vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10350__A1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] net922 vssd1
+ vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__and3_1
XANTENNA__09099__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14092__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08513_ net1070 net910 vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__and2_4
XFILLER_0_72_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ net548 _05686_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout256_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08444_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\] net726 _04684_
+ _04697_ _04647_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_92_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11850__A1 _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09859__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08763__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11470__B team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12058__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08375_ net1122 net961 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__and2_2
XFILLER_0_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout423_A _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10086__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13355__A1 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08271__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09594__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10814__B _06992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11198__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16474__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13107__B2 _03723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1407 net1412 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout420 net422 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
Xfanout431 _08023_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 _08021_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout453 _08018_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12521__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout464 net466 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_6
Xfanout475 net478 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_6
Xfanout486 _04556_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout497 _07810_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__dlymetal6s2s_1
X_09829_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\] net873 vssd1
+ vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12881__A3 _03589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ net3027 net284 net368 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14083__A2 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12771_ net2286 net198 net375 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XANTENNA__13291__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14510_ net1361 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
X_11722_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _07862_ vssd1 vssd1
+ vccd1 vccd1 _07863_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ net1266 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11841__B2 _07961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14441_ net1383 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
X_11653_ net2026 net1157 net567 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1
+ vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10604_ _06856_ _06858_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__or2_2
X_17160_ clknet_leaf_62_wb_clk_i _02720_ _01023_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14372_ net1326 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11584_ _04720_ _06847_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13323_ net119 net814 net807 net1746 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16111_ net1369 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] net715 _06782_ _06784_
+ _06787_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__a2111o_1
Xwire854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17091_ clknet_leaf_119_wb_clk_i _02651_ _00954_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16817__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire876 _04748_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16042_ net1405 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__inv_2
X_13254_ net602 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__inv_2
XANTENNA__13346__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\] net940
+ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__and3_1
X_12205_ net2763 net202 net441 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13185_ net2101 net1657 net828 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08222__B1 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ _06657_ _06658_ _06659_ _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12136_ net3240 net191 net447 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17993_ clknet_leaf_59_wb_clk_i _03542_ _01813_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11109__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13527__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12431__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12067_ _07841_ net494 _08012_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__and3_1
X_16944_ clknet_leaf_24_wb_clk_i _02504_ _00807_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09722__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ _07144_ _07278_ _07281_ _06970_ net545 vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__a221o_1
XANTENNA__08848__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16875_ clknet_leaf_46_wb_clk_i _02435_ _00738_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ net1179 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__inv_2
XANTENNA__10883__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15757_ net1214 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XANTENNA__13282__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ net1851 net606 net588 _03653_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a22o_1
XANTENNA__08828__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16139__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ net1374 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09679__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15688_ net1209 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17427_ clknet_leaf_50_wb_clk_i _02987_ _01290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__B _07553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14639_ net1364 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap855_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13585__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ net1688 net551 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1
+ vccd1 vccd1 _03535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18088__1462 vssd1 vssd1 vccd1 vccd1 _18088__1462/HI net1462 sky130_fd_sc_hd__conb_1
X_17358_ clknet_leaf_52_wb_clk_i _02918_ _01221_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10399__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08880__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16309_ clknet_leaf_112_wb_clk_i _01943_ _00177_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ net1063 team_01_WB.instance_to_wrap.cpu.f0.num\[17\] vssd1 vssd1 vccd1 vccd1
+ _04520_ sky130_fd_sc_hd__nand2_1
X_17289_ clknet_leaf_38_wb_clk_i _02849_ _01152_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12606__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17742__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09005__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10353__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08993_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] net886
+ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__and3_1
XANTENNA__17892__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12341__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__C_N _06992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout373_A _03571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] net655 _05862_ _05865_
+ _05872_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09545_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\] net651 _05792_ _05795_
+ _05806_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout540_A _06382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1282_A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13812__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16049__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13172__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] net644 net610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\]
+ _05732_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17272__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ net1142 net925 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14792__A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout805_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09886__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10528__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13576__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\] _04621_ vssd1 vssd1 vccd1 vccd1
+ _04622_ sky130_fd_sc_hd__and4_2
XFILLER_0_18_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ net2427 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12516__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] net751 _04651_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\]
+ _06564_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11339__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\] net625 _06491_ _06495_
+ _06505_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10263__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ _06442_ _06443_ _06444_ _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10562__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1207 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1218 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_2
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12251__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1240 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_4
X_14990_ net1231 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
Xfanout250 net253 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_2
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_4
Xfanout261 _07989_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
XANTENNA__13500__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1259 net1260 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_4
XANTENNA__13500__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 _07957_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
X_13941_ net1163 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[22\] sky130_fd_sc_hd__and3b_1
Xfanout283 _07920_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_1
Xfanout294 net297 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XFILLER_0_9_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16660_ clknet_leaf_104_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[14\]
+ _00523_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13872_ _04560_ _07680_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ net1298 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12823_ net3167 _07994_ net374 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
X_16591_ clknet_leaf_66_wb_clk_i _02219_ _00454_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13264__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15542_ net1260 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ net2366 net244 net381 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
XANTENNA__09499__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11705_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__and2_2
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ net2099 net263 net388 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ net1199 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_144_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11027__C1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17212_ clknet_leaf_16_wb_clk_i _02772_ _01075_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14424_ net1279 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
X_11636_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[8\] _07806_ vssd1 vssd1 vccd1
+ vccd1 _07833_ sky130_fd_sc_hd__and2_1
X_18192_ net1566 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
XANTENNA__09235__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__B _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17143_ clknet_leaf_12_wb_clk_i _02703_ _01006_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11567_ _07722_ _07734_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1
+ vccd1 _07793_ sky130_fd_sc_hd__a21o_1
X_14355_ net1655 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12426__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11330__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ net117 net811 net806 net1712 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
X_10518_ net971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] net956 vssd1
+ vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__and3_1
Xhold709 team_01_WB.instance_to_wrap.cpu.f0.num\[12\] vssd1 vssd1 vccd1 vccd1 net2325
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17074_ clknet_leaf_31_wb_clk_i _02634_ _00937_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14286_ _04193_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11498_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] _07721_ _07745_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\]
+ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13237_ _03721_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] net829 vssd1 vssd1
+ vccd1 vccd1 _02021_ sky130_fd_sc_hd__mux2_1
X_16025_ net1365 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\] net660 net642 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__a22o_1
XANTENNA__10002__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10173__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ net2713 net2501 net826 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09962__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12119_ net2195 net276 net453 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__mux2_1
XANTENNA__12161__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17976_ clknet_leaf_78_wb_clk_i _03525_ _01796_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13099_ net2135 net837 net357 _03719_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a22o_1
XANTENNA__10470__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1409 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net3025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16927_ clknet_leaf_1_wb_clk_i _02487_ _00790_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11502__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16858_ clknet_leaf_35_wb_clk_i _02418_ _00721_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10856__A2 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15809_ net1290 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16789_ clknet_leaf_8_wb_clk_i _02349_ _00652_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10069__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09330_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] net886
+ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10629__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\] net877 vssd1
+ vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08212_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__or4_1
XANTENNA__15501__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11018__C1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09192_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] net881
+ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ net1760 net552 net349 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1
+ vccd1 vccd1 _03552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11033__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12336__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout219_A _07925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08074_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 _04504_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_113_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1128_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A _03585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1 vccd1
+ net1630 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 _02122_ vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 net145 vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11195__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\] vssd1 vssd1 vccd1 vccd1 net1663
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold58 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\] vssd1 vssd1 vccd1 vccd1
+ net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] vssd1 vssd1 vccd1 vccd1
+ net1685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout755_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16662__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\] net856 vssd1
+ vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09459_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] net877
+ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08673__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13549__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ net3249 net204 net413 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08951__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] net1162 vssd1 vssd1 vccd1 vccd1
+ _07682_ sky130_fd_sc_hd__or2_2
XANTENNA__12246__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14140_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] _04242_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\]
+ _04291_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__a221o_1
XANTENNA__08976__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11352_ net339 net342 _05278_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10783__A1 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] net926 vssd1
+ vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14071_ net788 net787 _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__and3_4
XFILLER_0_46_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17168__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11283_ net541 _07408_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13022_ net1029 _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input51_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] net896 vssd1
+ vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__and3_1
XANTENNA__09782__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 net1008 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ clknet_leaf_88_wb_clk_i _03387_ _01651_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1012 _04484_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
X_10165_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] net883 vssd1
+ vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_2
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1045 net1046 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1
+ net1056 sky130_fd_sc_hd__clkbuf_4
X_17761_ clknet_leaf_89_wb_clk_i _03319_ _01582_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14973_ net1282 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
X_10096_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] net869 vssd1
+ vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__and3_1
Xfanout1067 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1
+ net1067 sky130_fd_sc_hd__clkbuf_4
Xfanout1078 net1080 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__dlymetal6s2s_1
X_18087__1461 vssd1 vssd1 vccd1 vccd1 _18087__1461/HI net1461 sky130_fd_sc_hd__conb_1
Xfanout1089 net1091 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_2
X_16712_ clknet_leaf_46_wb_clk_i _02272_ _00575_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13924_ net1166 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[5\] sky130_fd_sc_hd__and3b_1
X_17692_ clknet_leaf_82_wb_clk_i _03252_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16643_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[29\]
+ _00506_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11833__B _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13855_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] _04116_ net2434 vssd1 vssd1
+ vccd1 vccd1 _04136_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12806_ net2864 net224 net373 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16574_ clknet_leaf_142_wb_clk_i _02202_ _00437_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13786_ _04558_ _04084_ _04090_ net782 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o31a_1
X_10998_ net546 _07261_ _07079_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11799__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15525_ net1233 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XANTENNA__09022__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12737_ net2343 net289 net379 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XANTENNA__08664__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11263__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13540__S net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10168__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15456_ net1252 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
XANTENNA__09208__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12668_ net3197 net205 net389 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09957__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14201__A2 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14407_ net1309 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
X_18175_ net1549 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XANTENNA__12156__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ net497 _07824_ net2338 net839 vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o2bb2a_1
X_15387_ net1316 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XANTENNA__10465__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ net2177 net192 net395 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10223__B1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ clknet_leaf_141_wb_clk_i _02686_ _00989_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14338_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1
+ vccd1 _02260_ sky130_fd_sc_hd__clkbuf_1
Xhold506 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10774__A1 _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1 vccd1
+ net2133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11995__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold539 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ clknet_leaf_136_wb_clk_i _02617_ _00920_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\] _04239_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16008_ net1374 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_41_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15991__A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\] net752 net698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a22o_1
XANTENNA__14268__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1206 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08761_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] net936
+ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__and3_1
Xhold1228 team_01_WB.instance_to_wrap.cpu.K0.count\[1\] vssd1 vssd1 vccd1 vccd1 net2844
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ clknet_leaf_108_wb_clk_i net2856 _01779_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1239 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\] vssd1 vssd1 vccd1 vccd1
+ net2855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08692_ _04954_ _04955_ net580 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__mux2_1
XANTENNA__17930__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__A2 _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13779__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09447__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] net733 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\]
+ _05559_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a221o_1
XANTENNA__08655__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1078_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] net749 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09175_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\] net724 net721 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a22o_1
XANTENNA__12066__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout503_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04554_ vssd1 vssd1 vccd1 vccd1
+ _04555_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ team_01_WB.instance_to_wrap.cpu.f0.num\[29\] vssd1 vssd1 vccd1 vccd1 _04488_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1412_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout872_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14259__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08959_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\] net924
+ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11970_ net3257 net191 net467 vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__mux2_1
XANTENNA__09686__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10921_ net545 net531 _06953_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__and3_2
XFILLER_0_93_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11145__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ net541 _07115_ _07112_ _07111_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__o2bb2a_1
X_13640_ _07959_ _03972_ net187 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13571_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _05134_ _03902_ vssd1
+ vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a21oi_1
X_10783_ _05515_ _05448_ net508 vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15310_ net1229 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12522_ net2204 net317 net409 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16290_ clknet_leaf_98_wb_clk_i _01924_ _00158_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15241_ net1210 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
X_12453_ net2357 net266 net417 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10205__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11404_ net1155 _07662_ _07664_ _07666_ _07667_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__o311ai_2
XANTENNA__16558__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12384_ net2268 net276 net424 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
X_15172_ net1224 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XANTENNA__10756__A1 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17803__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18228__1589 vssd1 vssd1 vccd1 vccd1 _18228__1589/HI net1589 sky130_fd_sc_hd__conb_1
X_11335_ _06943_ _06945_ net322 _07588_ _07598_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__o41ai_1
X_14123_ _04153_ _04257_ _04259_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12704__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14054_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] _04218_ net565 vssd1
+ vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a21boi_1
X_11266_ _06954_ _07043_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__nand2_1
XANTENNA__10508__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08177__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\] net706 _06457_ _06462_
+ _06465_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a2111o_1
X_13005_ net2030 net248 net360 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11197_ _06347_ _06382_ _07459_ _07460_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17953__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__B2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17813_ clknet_leaf_68_wb_clk_i _03370_ _01634_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_10148_ _06402_ _06404_ _06408_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__or4_4
XFILLER_0_101_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17744_ clknet_leaf_105_wb_clk_i _03302_ _01565_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_10079_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] net740 net733 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__a22o_1
X_14956_ net1266 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XANTENNA__08856__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ net2683 net795 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[20\]
+ sky130_fd_sc_hd__and2_1
X_17675_ clknet_leaf_75_wb_clk_i _03235_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14887_ net1199 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
XANTENNA__10692__A0 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ clknet_leaf_105_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[12\]
+ _00489_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13838_ _04116_ _04126_ _04128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[9\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__09429__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16557_ clknet_leaf_23_wb_clk_i _02185_ _00420_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12433__A1 _07869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ net563 _04072_ _04075_ _04077_ _00020_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__a32o_1
XANTENNA__16147__A net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17333__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10444__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15508_ net1241 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16488_ clknet_leaf_106_wb_clk_i _02116_ _00351_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10995__A1 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10995__B2 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18227_ net602 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
X_15439_ net1248 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XANTENNA__10195__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09984__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18158_ net1532 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_0_68_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17483__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10747__A1 _07010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold314 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ clknet_leaf_8_wb_clk_i _02669_ _00972_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold325 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ net1463 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12614__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13937__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold336 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\] vssd1 vssd1 vccd1 vccd1
+ net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_01_WB.instance_to_wrap.cpu.c0.count\[14\] vssd1 vssd1 vccd1 vccd1 net1963
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\] net922 vssd1
+ vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__and3_1
XANTENNA__11738__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_2
XFILLER_0_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout816 _03740_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
Xfanout827 net832 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
X_09862_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\] net747 net722 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__a22o_1
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10361__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout849 _04769_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08573__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1003 team_01_WB.instance_to_wrap.cpu.f0.num\[4\] vssd1 vssd1 vccd1 vccd1 net2619
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08813_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\] net920
+ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and3_1
Xhold1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] net750 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a22o_1
Xhold1025 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1036 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout286_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15226__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1058 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _04999_ _05000_ _05002_ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1069 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\] vssd1 vssd1 vccd1 vccd1
+ net2685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\] net661 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\]
+ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout453_A _08018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1195_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08628__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A2 _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__B net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1362_A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13180__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10435__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08274__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09597__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17826__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09227_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] net924
+ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18086__1460 vssd1 vssd1 vccd1 vccd1 _18086__1460/HI net1460 sky130_fd_sc_hd__conb_1
XANTENNA__09894__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09158_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] net937
+ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08109_ _04475_ team_01_WB.instance_to_wrap.cpu.f0.num\[10\] _04498_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a221o_1
XANTENNA__12524__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09089_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\] net921
+ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__and3_1
XANTENNA__16850__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17976__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11120_ net333 _07382_ _07383_ _06175_ _06141_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11648__B _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _07045_ _07051_ net514 vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__mux2_1
Xhold892 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\] vssd1 vssd1 vccd1 vccd1
+ net2508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10271__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] net751 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\]
+ _06249_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__a221o_1
XANTENNA__17206__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15136__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ net1357 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
X_15790_ net1215 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1570 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3186 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09134__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1324 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
Xhold1581 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__B _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1592 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3208 sky130_fd_sc_hd__dlygate4sd3_1
X_11953_ net2758 net272 net471 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16230__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10904_ net514 _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__nand2_1
X_17460_ clknet_leaf_6_wb_clk_i _03020_ _01323_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14672_ net1402 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\] net678 net779 vssd1 vssd1
+ vccd1 vccd1 _07997_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16411_ clknet_leaf_100_wb_clk_i net2384 _00274_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13623_ net969 _03958_ _03954_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o21ai_1
X_17391_ clknet_leaf_53_wb_clk_i _02951_ _01254_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08619__B1 _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10835_ _07085_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10426__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16342_ clknet_leaf_63_wb_clk_i net1669 _00210_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08095__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13554_ net767 _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08095__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10766_ _06071_ _05852_ net504 vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__mux2_1
XANTENNA__09831__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12505_ net3246 net232 net408 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
X_16273_ clknet_leaf_66_wb_clk_i _01910_ _00141_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09300__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13485_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _05380_ _05449_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a22o_1
X_10697_ _05448_ _05378_ net502 vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ net107 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
X_15224_ net1257 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
X_12436_ net3195 net241 net417 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11839__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ net1186 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12434__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12367_ net2764 net194 net425 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ net792 _04228_ _04243_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__and3_4
XFILLER_0_107_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _06721_ _07124_ _06720_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__a21bo_1
X_12298_ net1926 net214 net434 vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
X_15086_ net1228 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14037_ net565 _04208_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__and2_1
X_11249_ net324 _07512_ _06920_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__or3b_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11154__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08570__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15988_ net1381 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__inv_2
X_17727_ clknet_leaf_96_wb_clk_i _03285_ _01548_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14939_ net1317 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ net772 net766 net681 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__or3_1
X_17658_ clknet_leaf_36_wb_clk_i _03218_ _01521_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08883__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16723__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16609_ clknet_leaf_111_wb_clk_i _02237_ _00472_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17849__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08391_ net1153 net1151 net1149 net1148 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and4b_4
XANTENNA__12609__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17589_ clknet_leaf_26_wb_clk_i _03149_ _01452_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10918__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10417__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12957__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16873__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09012_ _05272_ _05274_ _05275_ _05245_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o31a_4
XANTENNA__10356__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09035__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11749__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\] vssd1 vssd1 vccd1 vccd1
+ net1727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A _07906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 net1738
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold133 net98 vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\] vssd1 vssd1 vccd1 vccd1
+ net1760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17229__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__B net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\] vssd1 vssd1 vccd1 vccd1
+ net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold177 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_2
Xhold199 net108 vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _06071_ _06108_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__xor2_4
XFILLER_0_10_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout613 _04775_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_4
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout635 _04761_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_6
XANTENNA__10091__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1208_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 _04751_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_8
Xfanout657 _04740_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_8
X_09845_ _06071_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nor2_1
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_8
XANTENNA__09880__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__B2 _03598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout668_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08561__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14095__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _05852_ _05889_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\] net638 net610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09889__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] net686 _04910_
+ _04913_ _04917_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_55_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12519__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ _04828_ _04851_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12948__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _06456_ _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13070__A1 _05480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\] net662 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\]
+ _06814_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__a221o_1
XANTENNA__09120__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _06724_ _06743_ _06744_ _06745_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__or4_1
X_13270_ net88 net816 net600 net2467 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ net2641 net268 net442 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12254__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A2 _06450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12152_ net2611 net275 net448 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__mux2_1
XANTENNA__09129__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08033__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11899__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _06869_ _07351_ _07355_ _07363_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12083_ net2559 net280 net456 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__mux2_1
X_16960_ clknet_leaf_142_wb_clk_i _02520_ _00823_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15911_ net1383 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__inv_2
X_11034_ _05069_ net340 _07297_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16891_ clknet_leaf_32_wb_clk_i _02451_ _00754_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09790__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08552__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ net1266 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14086__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16746__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ net1278 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12636__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ team_01_WB.instance_to_wrap.a1.ADR_I\[0\] net604 net586 _03664_ vssd1 vssd1
+ vccd1 vccd1 _02208_ sky130_fd_sc_hd__a22o_1
X_17512_ clknet_leaf_62_wb_clk_i _03072_ _01375_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ net1320 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11936_ net2663 net206 net473 vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17443_ clknet_leaf_119_wb_clk_i _03003_ _01306_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14655_ net1364 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12429__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\] net677 net779 vssd1 vssd1
+ vccd1 vccd1 _07983_ sky130_fd_sc_hd__o21a_1
XANTENNA__10738__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16896__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ net772 _07520_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10818_ net346 _07024_ _07026_ _07081_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a211o_1
X_17374_ clknet_leaf_12_wb_clk_i _02934_ _01237_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14586_ net1411 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _07857_ vssd1 vssd1
+ vccd1 vccd1 _07926_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16325_ clknet_leaf_64_wb_clk_i net1699 _00193_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13537_ _03861_ _03863_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__xor2_1
X_10749_ _06141_ _06071_ net507 vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16256_ clknet_leaf_69_wb_clk_i _01893_ _00124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13468_ _03816_ _03819_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09965__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15207_ net1180 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
X_12419_ net2606 net270 net419 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
XANTENNA__12164__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16187_ clknet_leaf_86_wb_clk_i _01854_ _00055_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10473__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10178__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _04850_ vssd1 vssd1
+ vccd1 vccd1 _03752_ sky130_fd_sc_hd__nand2_1
X_15138_ net1263 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08791__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15069_ net1281 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XANTENNA__17521__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08878__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12875__B2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] net963
+ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__and3_1
XANTENNA__10350__A2 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] net943 vssd1
+ vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08512_ net1081 net845 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_2
X_09492_ _05688_ _05755_ _05689_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09502__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08443_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] net717 _04686_ _04689_
+ _04692_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12339__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout249_A _07953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ net1148 net1150 net1153 net1152 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_110_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17051__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12074__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16619__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1325_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11198__B _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13694__A team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08782__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1408 net1412 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__buf_2
Xfanout410 _03562_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 _08023_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16769__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 _08020_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout454 _08018_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_A _04644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_8
Xfanout476 net478 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] net879 vssd1
+ vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__and3_1
Xfanout498 net500 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
X_09759_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] net645 _05995_
+ _05998_ _06004_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13633__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ net3231 net286 net375 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13291__B2 team_01_WB.instance_to_wrap.a1.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_115_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11721_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ _07861_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__and3_1
XANTENNA__12249__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14440_ net1382 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11652_ net1969 net1157 net567 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1
+ vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09247__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13942__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14240__B1 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10603_ _06858_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14371_ net1326 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11583_ _04720_ _06847_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__and2_2
XFILLER_0_92_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16110_ net1356 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13322_ net2258 net813 net807 net2156 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a22o_1
X_10534_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] net720 net717 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__a221o_1
X_17090_ clknet_leaf_144_wb_clk_i _02650_ _00953_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09785__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16041_ net1365 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__inv_2
XANTENNA__13346__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13253_ _03732_ _03733_ _03734_ _03737_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__or4_1
XFILLER_0_122_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10465_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\] net931
+ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17544__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ net2574 net239 net441 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_1
X_13184_ net2827 net2805 net826 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
X_10396_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\] net623 _04773_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\] _06646_ vssd1 vssd1 vccd1
+ vccd1 _06660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ net2554 net196 net449 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__mux2_1
XANTENNA__08773__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17992_ clknet_leaf_64_wb_clk_i _03541_ _01812_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12712__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16943_ clknet_leaf_18_wb_clk_i _02503_ _00806_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12066_ net2824 net210 net462 vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__B _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _07279_ _07280_ net528 vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__mux2_1
X_16874_ clknet_leaf_47_wb_clk_i _02434_ _00737_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15825_ net1195 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__inv_2
XANTENNA__09025__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18065__1439 vssd1 vssd1 vccd1 vccd1 _18065__1439/HI net1439 sky130_fd_sc_hd__conb_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15756_ net1286 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
X_12968_ net365 _03651_ _03652_ net1055 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09322__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ net1371 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11919_ net3019 net246 net475 vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12159__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15687_ net1195 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] net1056 net366 _03602_
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17426_ clknet_leaf_39_wb_clk_i _02986_ _01289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14638_ net1375 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XANTENNA__17074__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14231__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17357_ clknet_leaf_19_wb_clk_i _02917_ _01220_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14569_ net1334 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ clknet_leaf_111_wb_clk_i _01942_ _00176_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08090_ net1063 team_01_WB.instance_to_wrap.cpu.f0.num\[17\] vssd1 vssd1 vccd1 vccd1
+ _04519_ sky130_fd_sc_hd__or2_1
X_17288_ clknet_leaf_45_wb_clk_i _02848_ _01151_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15994__A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16239_ clknet_leaf_79_wb_clk_i _00019_ _00107_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13337__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09992__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16911__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12622__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\] net851 vssd1
+ vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08401__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08516__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09613_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\] net896 vssd1
+ vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout366_A _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\] net660 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a22o_1
XANTENNA__09477__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17417__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09232__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12069__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11823__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] net655 _05723_
+ _05731_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout533_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1275_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08426_ net1142 _04677_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14222__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ net1156 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout700_A _04685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11587__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08282__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08288_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10250_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\] net631 _06497_ _06502_
+ _06507_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10181_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] net610 _06421_ _06428_
+ _06437_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12532__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_4
XANTENNA__10562__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1216 net1218 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_4
XANTENNA__08949__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1227 net1236 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
Xfanout1238 net1240 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_4
Xfanout1249 net1268 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_2
Xfanout251 net253 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xfanout262 net265 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_2
X_13940_ net1164 net1057 net1665 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[21\]
+ sky130_fd_sc_hd__and3b_1
Xfanout273 _07957_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
Xfanout284 _07920_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_2
Xfanout295 net297 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09180__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ team_01_WB.instance_to_wrap.cpu.f0.state\[8\] _04566_ _04617_ net3078 vssd1
+ vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15610_ net1305 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
X_12822_ net3059 net260 net373 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16590_ clknet_leaf_79_wb_clk_i _02218_ _00453_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17097__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15541_ net1176 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12753_ net2073 net316 net382 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11704_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__and2b_1
X_15472_ net1250 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
X_12684_ net2264 net269 net389 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__mux2_1
XANTENNA__08981__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08691__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ clknet_leaf_39_wb_clk_i _02771_ _01074_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ net1280 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11635_ net1998 net840 _07808_ _07832_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__o22a_1
X_18191_ net1565 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
XANTENNA__12707__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17142_ clknet_leaf_32_wb_clk_i _02702_ _01005_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14354_ net3187 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _04480_ _07731_ _07769_ _07792_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16934__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13319__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13305_ net118 net809 net804 net1751 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a22o_1
X_17073_ clknet_leaf_21_wb_clk_i _02633_ _00936_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10517_ net971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] net948 vssd1
+ vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and3_1
X_14285_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _04436_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ _07724_ _07734_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_113_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16024_ net1377 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13236_ _03720_ net2158 net819 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_1
X_10448_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\] net656 net610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\]
+ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13167_ net1771 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\] net830 vssd1 vssd1
+ vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
XANTENNA__10751__A _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12442__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10379_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] net759 _06641_ _06642_
+ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10553__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ net1970 net215 net451 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__mux2_1
X_17975_ clknet_leaf_70_wb_clk_i _03524_ _01795_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13098_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\] _06106_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16926_ clknet_leaf_12_wb_clk_i _02486_ _00789_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ net2924 net251 net459 vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11502__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16857_ clknet_leaf_18_wb_clk_i _02417_ _00720_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11582__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15808_ net1272 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
X_16788_ clknet_leaf_6_wb_clk_i _02348_ _00651_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08594__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739_ net1299 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_18029__1423 vssd1 vssd1 vccd1 vccd1 _18029__1423/HI net1423 sky130_fd_sc_hd__conb_1
XFILLER_0_133_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10198__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap965_A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16464__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09987__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\] net842
+ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14204__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04574_ vssd1 vssd1 vccd1 vccd1
+ _04606_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09191_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] net871
+ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__and3_1
X_17409_ clknet_leaf_136_wb_clk_i _02969_ _01272_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12617__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08142_ _04566_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10645__B _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08073_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] vssd1 vssd1 vccd1 vccd1 _04503_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10792__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08737__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09227__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__B _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ net712 _05231_ _05235_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__or4_4
XFILLER_0_23_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout483_A _07702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\] vssd1 vssd1 vccd1 vccd1 net1631
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 team_01_WB.instance_to_wrap.a1.ADR_I\[8\] vssd1 vssd1 vccd1 vccd1 net1642
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\] vssd1 vssd1 vccd1 vccd1
+ net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold48 _02119_ vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] vssd1 vssd1 vccd1 vccd1
+ net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1392_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11492__A _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08277__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09527_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] _04772_ vssd1
+ vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12100__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09897__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] net882 vssd1
+ vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16957__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13549__A2 _07653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08409_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] net954 vssd1
+ vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__and3_1
XANTENNA__12527__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _05243_ net577 vssd1 vssd1
+ vccd1 vccd1 _05653_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11420_ net785 _07680_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ net538 _07475_ _07471_ _07002_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] net963 vssd1
+ vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__and3_1
X_14070_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nor2_2
X_18064__1438 vssd1 vssd1 vccd1 vccd1 _18064__1438/HI net1438 sky130_fd_sc_hd__conb_1
XFILLER_0_123_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _07179_ _07184_ net539 vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13021_ _04795_ net571 _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08728__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] net892 vssd1
+ vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12262__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10535__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\] net869 vssd1
+ vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__and3_1
Xfanout1002 net1004 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09137__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__A team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1024 _04484_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1 vccd1 net1046
+ sky130_fd_sc_hd__clkbuf_4
X_14972_ net1234 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
X_10095_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] net853 vssd1
+ vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17760_ clknet_leaf_89_wb_clk_i _03318_ _01581_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1057 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1057 sky130_fd_sc_hd__clkbuf_2
Xfanout1068 net1071 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_2
XANTENNA__13485__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1079 net1080 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XANTENNA__13485__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16711_ clknet_leaf_121_wb_clk_i _02271_ _00574_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13923_ net1165 net1059 net3073 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[4\]
+ sky130_fd_sc_hd__and3b_1
X_17691_ clknet_leaf_84_wb_clk_i _03251_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16642_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[28\]
+ _00505_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13854_ _04115_ _04135_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[8\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13237__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17732__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ net2333 net229 net371 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16573_ clknet_leaf_136_wb_clk_i _02201_ _00436_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09303__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13785_ _04473_ _07776_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__and2_1
X_10997_ net534 _07260_ _07250_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_1389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15524_ net1269 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XANTENNA__15602__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12736_ net2365 net232 net380 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17882__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09600__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15455_ net1295 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12437__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ net2754 net238 net387 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ net1308 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
X_18174_ net1548 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XFILLER_0_5_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11618_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[17\] net573 vssd1 vssd1 vccd1
+ vccd1 _07824_ sky130_fd_sc_hd__nand2_1
X_15386_ net1259 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
X_12598_ net2239 net194 net395 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ clknet_leaf_133_wb_clk_i _02685_ _00988_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10223__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14337_ net1966 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11549_ net483 _07781_ net319 vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__a21o_1
XANTENNA__17112__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold507 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold518 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold529 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ clknet_leaf_142_wb_clk_i _02616_ _00919_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\] _04229_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\]
+ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16007_ net1368 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__inv_2
X_13219_ net2383 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\] net825 vssd1 vssd1
+ vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
XANTENNA__12172__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14199_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\] _04252_ _04278_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\]
+ _04354_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1207 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08760_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] net944 vssd1
+ vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__and3_1
X_17958_ clknet_leaf_104_wb_clk_i _03508_ _01778_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ sky130_fd_sc_hd__dfstp_1
Xhold1218 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_81_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1229 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08886__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09144__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16909_ clknet_leaf_19_wb_clk_i _02469_ _00772_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_08691_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net763 net590 vssd1 vssd1
+ vccd1 vccd1 _04955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17889_ clknet_leaf_109_wb_clk_i _03439_ _01709_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13779__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09312_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] net741 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\]
+ _05554_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a221o_1
XANTENNA__10359__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] net729 net725 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\]
+ _05495_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a221o_1
XANTENNA__12347__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout231_A _07897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _05434_ _05435_ _05436_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ _04551_ _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__nor2_1
XANTENNA__11411__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1140_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09080__B2 _05343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ net1156 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__inv_2
XANTENNA__09883__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13178__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout698_A _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12082__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1405_A net1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12911__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14798__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\] net922
+ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__and3_1
XANTENNA__12810__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08889_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\] net754 net746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\]
+ _05142_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a221o_1
X_10920_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10150__B1 _06412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ _07113_ _07114_ net529 vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09123__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10269__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ net966 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _03912_ _03913_
+ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10782_ _07044_ _07045_ net514 vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10453__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12521_ net2194 net303 net409 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
XANTENNA__11650__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12257__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17135__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10566__A _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15240_ net1208 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12452_ net2988 net270 net415 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
XANTENNA__08036__A team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11403_ _04486_ _07023_ _07665_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15171_ net1220 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12383_ net2244 net217 net423 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XANTENNA__11953__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14122_ _04265_ _04271_ _04277_ _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__or4_1
X_11334_ _07004_ _07546_ _07589_ _07079_ _07597_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_65_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11397__A _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ _04218_ net565 _04217_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__and3b_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18028__1422 vssd1 vssd1 vccd1 vccd1 _18028__1422/HI net1422 sky130_fd_sc_hd__conb_1
X_11265_ net544 _07528_ _07527_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13004_ net2027 net277 net362 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
X_10216_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] net753 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__a22o_1
X_11196_ _06384_ _06983_ _06985_ net536 net331 vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11181__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17812_ clknet_leaf_68_wb_clk_i _03369_ _01633_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_10147_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\] net723 net714 _06409_
+ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12720__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14955_ net1205 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
X_17743_ clknet_leaf_104_wb_clk_i _03301_ _01564_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_10078_ _06338_ _06339_ _06340_ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__or4_1
XFILLER_0_136_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] net795 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[19\] sky130_fd_sc_hd__and2_1
X_17674_ clknet_leaf_73_wb_clk_i _03234_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14886_ net1314 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13837_ team_01_WB.instance_to_wrap.cpu.c0.count\[9\] _04115_ vssd1 vssd1 vccd1 vccd1
+ _04128_ sky130_fd_sc_hd__or2_1
XANTENNA__10692__A1 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16625_ clknet_leaf_96_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[11\]
+ _00488_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12969__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16556_ clknet_leaf_30_wb_clk_i _02184_ _00419_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13768_ _07713_ _04076_ net784 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18179__1553 vssd1 vssd1 vccd1 vccd1 _18179__1553/HI net1553 sky130_fd_sc_hd__conb_1
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09330__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12719_ net2464 net305 net383 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
X_15507_ net1189 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16487_ clknet_leaf_76_wb_clk_i _02115_ _00350_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13699_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _04020_ vssd1 vssd1 vccd1 vccd1
+ _04021_ sky130_fd_sc_hd__or2_1
X_15438_ net1231 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
X_18226_ net602 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16502__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18157_ net1531 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
X_15369_ net1210 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17108_ clknet_leaf_6_wb_clk_i _02668_ _00971_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold304 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ net1462 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_106_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold315 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold326 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 team_01_WB.instance_to_wrap.a1.ADR_I\[26\] vssd1 vssd1 vccd1 vccd1 net1953
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[3\] vssd1 vssd1 vccd1 vccd1 net1964
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09930_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] net942 vssd1
+ vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__and3_1
X_17039_ clknet_leaf_54_wb_clk_i _02599_ _00902_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold359 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17778__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout806 net807 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_2
X_09861_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\] net915 vssd1
+ vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__and3_1
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
Xfanout828 net832 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_4
Xfanout839 team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1
+ net839 sky130_fd_sc_hd__buf_2
X_08812_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] _04644_
+ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__and3_1
Xhold1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] net740 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a22o_1
Xhold1015 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 net2631
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14411__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17008__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1026 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _05003_ _05004_ _05005_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or4_1
Xhold1048 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08674_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[28\] net664 net635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18063__1437 vssd1 vssd1 vccd1 vccd1 _18063__1437/HI net1437 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout446_A _08020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1188_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12077__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout613_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09226_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\] net936 vssd1
+ vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14177__A2 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16182__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13697__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\] net913
+ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12805__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08108_ _04472_ team_01_WB.instance_to_wrap.cpu.f0.num\[15\] _04498_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08800__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ net1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] net918
+ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08039_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 _04470_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_13_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold860 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold871 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold882 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _06833_ net340 net338 _06830_ _07313_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__o221a_1
Xhold893 _03437_ vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09118__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12360__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__B1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10001_ _06262_ _06263_ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12540__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10371__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09108__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1560 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\] vssd1 vssd1 vccd1 vccd1
+ net3176 sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ net1319 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
Xhold1571 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ net3172 net246 net471 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux2_1
Xhold1582 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3209 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _04828_ _04883_ net498 vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__mux2_1
X_14671_ net1364 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11883_ net678 _07478_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16410_ clknet_leaf_102_wb_clk_i net2569 _00273_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15152__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13622_ _07535_ _03957_ net770 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17390_ clknet_leaf_55_wb_clk_i _02950_ _01253_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08619__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10834_ _07091_ _07097_ net539 vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13612__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09788__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16341_ clknet_leaf_63_wb_clk_i net1759 _00209_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13553_ _07898_ _03898_ net185 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10765_ _07027_ _07028_ net519 vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12504_ net3154 net236 net407 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
X_16272_ clknet_leaf_69_wb_clk_i _01909_ _00140_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13484_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _05244_ _05310_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__o211a_1
X_10696_ _06956_ _06959_ net514 vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18011_ clknet_leaf_79_wb_clk_i _03560_ _01825_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15223_ net1243 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ net3131 net207 net417 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
XANTENNA__09044__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12715__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11387__C1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13400__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ net1178 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XANTENNA__17920__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12366_ _07846_ _08011_ net488 vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14105_ net793 _04226_ _04241_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__and3_4
XFILLER_0_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ _07572_ _07579_ _07580_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__and3_1
X_15085_ net1212 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12297_ net2835 net291 net432 vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XANTENNA__10462__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] _04207_ vssd1 vssd1 vccd1
+ vccd1 _04208_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09347__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11248_ _05485_ _06919_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__nor2_1
XANTENNA__09028__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08555__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15327__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _06455_ _06594_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10362__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15987_ net1384 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11066__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17726_ clknet_leaf_96_wb_clk_i _03284_ _01547_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10114__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14938_ net1265 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11862__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17657_ clknet_leaf_125_wb_clk_i _03217_ _01520_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14869_ net1343 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ clknet_leaf_111_wb_clk_i _02236_ _00471_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_08390_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\] net945 vssd1
+ vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__and3_1
XANTENNA__09807__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17588_ clknet_leaf_4_wb_clk_i _03148_ _01451_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_16539_ clknet_leaf_61_wb_clk_i _02167_ _00402_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09995__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14159__A2 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09011_ _05264_ _05265_ _05266_ _05267_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18209_ net1583 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
XANTENNA__12625__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14406__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 net1717
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11749__B _07585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\] vssd1 vssd1 vccd1 vccd1
+ net1728 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold123 _01982_ vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 _02013_ vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold145 net139 vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _02091_ vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\] vssd1 vssd1 vccd1 vccd1
+ net1794 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _06110_ _06176_ _06109_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__a21o_1
Xfanout603 net179 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_125_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold189 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] vssd1 vssd1 vccd1 vccd1
+ net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _04774_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_6
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout625 _04767_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_8
XFILLER_0_61_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout396_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout636 _04761_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12360__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout647 _04751_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_4
X_09844_ net581 _06105_ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__a21oi_4
Xfanout658 _04739_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout669 _04730_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_4
XANTENNA__12893__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ _05852_ _05889_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13980__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\] net618 net609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16548__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09510__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _04914_ _04918_ _04919_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout730_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08285__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ _04828_ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__and2_1
X_18027__1421 vssd1 vssd1 vccd1 vccd1 _18027__1421/HI net1421 sky130_fd_sc_hd__conb_1
XFILLER_0_14_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16218__D team_01_WB.instance_to_wrap.cpu.c0.next_atmax vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16698__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15700__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17943__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] net616 net610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__a22o_1
X_09209_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\] net625 _05456_ _05463_
+ _05465_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13358__B1 _03747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10481_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\] net719 _06732_
+ _06735_ _06737_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12535__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ net2818 net271 net439 vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09577__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08785__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ net2137 net218 net447 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__mux2_1
XANTENNA__10282__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ net547 _07365_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ net2408 net250 net457 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__mux2_1
Xhold690 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18178__1552 vssd1 vssd1 vccd1 vccd1 _18178__1552/HI net1552 sky130_fd_sc_hd__conb_1
X_11033_ _05068_ net338 net332 _05066_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__o221a_1
X_15910_ net1341 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__inv_2
XANTENNA__12270__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890_ clknet_leaf_34_wb_clk_i _02450_ _00753_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11394__B _07551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ net1313 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_138_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ net1278 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
X_12984_ _07121_ _03662_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] net1053
+ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__a2bb2o_1
Xhold1390 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\] vssd1 vssd1 vccd1 vccd1
+ net3006 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17511_ clknet_leaf_131_wb_clk_i _03071_ _01374_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14723_ net1320 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11935_ net2954 net190 net471 vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17442_ clknet_leaf_142_wb_clk_i _03002_ _01305_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14654_ net1378 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
X_11866_ net677 _07396_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__nand2_1
XANTENNA__10738__B _06995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ _07936_ _03942_ net186 vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__mux2_1
XANTENNA__13114__B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817_ _07004_ _07043_ _07077_ _07079_ _07068_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__a221o_1
XANTENNA__10951__A2_N net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14585_ net1411 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
X_17373_ clknet_leaf_127_wb_clk_i _02933_ _01236_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11797_ net2961 net220 net480 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16324_ clknet_leaf_76_wb_clk_i _01958_ _00192_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
X_13536_ net185 _07885_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor2_1
X_10748_ _06277_ _06211_ net507 vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13349__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16255_ clknet_leaf_69_wb_clk_i _01892_ _00123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _05719_ vssd1 vssd1
+ vccd1 vccd1 _03820_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10679_ _06935_ _06941_ _04959_ _06840_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15206_ net1271 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12418_ net3243 net247 net420 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XANTENNA__11569__B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16186_ clknet_leaf_97_wb_clk_i net840 _00054_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13398_ net2602 net327 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12572__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15137_ net1291 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12349_ net2150 net216 net490 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
X_18062__1436 vssd1 vssd1 vccd1 vccd1 _18062__1436/HI net1436 sky130_fd_sc_hd__conb_1
XFILLER_0_26_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15068_ net1280 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08528__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__or4b_1
XANTENNA__12180__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12875__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09055__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10886__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14896__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09560_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08511_ net994 net850 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__and2_2
X_17709_ clknet_leaf_109_wb_clk_i _03269_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09491_ _05718_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16840__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08442_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\] net721 net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10648__B _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11835__A1_N net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08373_ _04624_ _04635_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16990__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12355__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11479__B _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16220__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09891__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _03564_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_4
Xfanout1409 net1410 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__buf_4
XANTENNA__08519__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 _03561_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_6
Xfanout422 _08028_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13186__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout778_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 _08023_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout444 _08020_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_4
XANTENNA__12866__A2 _07834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 net458 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16370__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 _08014_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout477 net478 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_8
X_09827_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\] net865 vssd1
+ vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout488 _08026_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout945_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] net624 _06021_ net671
+ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a211o_1
XANTENNA__13815__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08709_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] net924 vssd1
+ vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11826__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09689_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\] net649 _05931_ _05947_
+ net672 vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__a2111o_1
X_11720_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _07860_ vssd1 vssd1
+ vccd1 vccd1 _07861_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11651_ net2147 net1157 net567 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1
+ vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a22o_1
XANTENNA__09131__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__B_N _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ _06863_ _06865_ _06860_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__or3b_2
X_14370_ net1326 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
XANTENNA__09798__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ net1161 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\] vssd1 vssd1 vccd1
+ vccd1 team_01_WB.instance_to_wrap.cpu.DM0.next_enable sky130_fd_sc_hd__and2_1
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ net133 net813 net807 net1964 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10533_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] net748 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12265__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ net1374 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13252_ net63 net62 _03735_ _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input74_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] net723 net690 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__a22o_1
Xwire889 net890 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08044__A team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ net2766 net207 net441 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ net2183 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\] net830 vssd1 vssd1
+ vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
X_10395_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\] net639 net608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\]
+ _06645_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ net495 _07845_ _08017_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__and3_4
XFILLER_0_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09970__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16713__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17991_ clknet_leaf_59_wb_clk_i _03540_ _01811_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ net2313 net291 net461 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux2_1
X_16942_ clknet_leaf_52_wb_clk_i _02502_ _00805_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10317__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11016_ _07028_ _07047_ net516 vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__mux2_1
XANTENNA__09722__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16873_ clknet_leaf_41_wb_clk_i _02433_ _00736_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11004__A2_N net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15605__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ net1253 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17989__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12967_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1
+ vccd1 _03652_ sky130_fd_sc_hd__or2_1
X_15755_ net1204 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13282__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ net1406 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
X_11918_ net2354 net274 net476 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15686_ net1271 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
X_12898_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] _07324_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17425_ clknet_leaf_22_wb_clk_i _02985_ _01288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14637_ net1369 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
X_11849_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _07851_ vssd1 vssd1 vccd1
+ vccd1 _07968_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ clknet_leaf_44_wb_clk_i _02916_ _01219_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14568_ net1334 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08880__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16307_ clknet_leaf_112_wb_clk_i _01941_ _00175_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16243__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12175__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] _03871_ net1067 vssd1
+ vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14499_ net1362 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17287_ clknet_leaf_120_wb_clk_i _02847_ _01150_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16238_ clknet_leaf_79_wb_clk_i _00018_ _00106_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16169_ clknet_leaf_57_wb_clk_i _01837_ _00037_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10556__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16393__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] net845
+ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18026__1420 vssd1 vssd1 vccd1 vccd1 _18026__1420/HI net1420 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\] net885 vssd1
+ vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09543_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] net885 vssd1
+ vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout261_A _07989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09474_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\] net842
+ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[31\] net941
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1170_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10097__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11036__A1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15250__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1268_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\] net3116 net1042 vssd1 vssd1
+ vccd1 vccd1 _03391_ sky130_fd_sc_hd__mux2_1
X_18177__1551 vssd1 vssd1 vccd1 vccd1 _18177__1551/HI net1551 sky130_fd_sc_hd__conb_1
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09886__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12085__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\]
+ net1044 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16736__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12813__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10547__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\] _04777_ _06417_
+ _06431_ _06434_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1206 net1207 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_4
Xfanout1217 net1218 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_2
Xfanout1228 net1235 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_4
Xfanout230 _07897_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout241 _07884_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_121_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_2
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_2
Xfanout263 net265 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
Xfanout274 _07948_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09126__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout285 _07920_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04555_ _04567_ _04141_ vssd1
+ vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12821_ net2842 net300 net374 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__mux2_1
XANTENNA__13264__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ net2903 net305 net380 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
X_15540_ net1237 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
XANTENNA__11391__C _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08039__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11703_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] _07835_ _07840_ vssd1 vssd1
+ vccd1 vccd1 _07844_ sky130_fd_sc_hd__and3_1
X_15471_ net1247 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XANTENNA__16266__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12683_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\] net270 net387 vssd1
+ vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08981__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ net1280 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
X_17210_ clknet_leaf_34_wb_clk_i _02770_ _01073_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15160__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17511__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[9\] _07806_ vssd1 vssd1 vccd1
+ vccd1 _07832_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18190_ net1564 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12775__A1 _07925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11122__S1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14353_ net1656 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17141_ clknet_leaf_26_wb_clk_i _02701_ _01004_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11565_ net320 _07791_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1
+ vccd1 _07792_ sky130_fd_sc_hd__o21a_1
XANTENNA__08443__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13304_ net120 net808 net803 net1971 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17072_ clknet_leaf_23_wb_clk_i _02632_ _00935_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10516_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\] net961
+ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10250__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14284_ _04201_ _04435_ net1367 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a21oi_1
X_11496_ _07742_ _07744_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1
+ vccd1 _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17661__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13235_ _03719_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] net831 vssd1 vssd1
+ vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16023_ net1376 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10447_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] net653 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12723__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10002__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09943__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10378_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12117_ net2001 net281 net453 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__mux2_1
XANTENNA__11750__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17974_ clknet_leaf_72_wb_clk_i _03523_ _01794_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13097_ net354 _03717_ _03718_ net835 net2962 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a32o_1
XANTENNA__10470__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ net2263 net255 net461 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
X_16925_ clknet_leaf_127_wb_clk_i _02485_ _00788_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12959__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16856_ clknet_leaf_26_wb_clk_i _02416_ _00719_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09333__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15807_ net1294 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16787_ clknet_leaf_47_wb_clk_i _02347_ _00650_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13999_ _04169_ _03553_ _04183_ _03558_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__a31o_1
XANTENNA__10069__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15738_ net1307 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15669_ net1177 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17191__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11802__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _04568_ _04604_ _04605_ net553 net1653 vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17408_ clknet_leaf_140_wb_clk_i _02968_ _01271_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_09190_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] net851
+ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16759__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08141_ team_01_WB.instance_to_wrap.cpu.f0.state\[7\] net553 vssd1 vssd1 vccd1 vccd1
+ _04568_ sky130_fd_sc_hd__nor2_2
X_17339_ clknet_leaf_37_wb_clk_i _02899_ _01202_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08434__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] vssd1 vssd1 vccd1 vccd1 _04502_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13715__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12518__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12633__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14414__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08198__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09508__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08412__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10661__B _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ _05225_ _05226_ _05236_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout1016_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 _03410_ vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold27 _01991_ vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14140__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13932__A_N net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\] vssd1 vssd1 vccd1 vccd1
+ net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 net1665
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15245__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10701__A0 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout643_A _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1385_A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\] net910 vssd1
+ vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__and3_1
XANTENNA__17534__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] net666 vssd1 vssd1
+ vccd1 vccd1 _05721_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout810_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12808__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ net984 net954 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and2_4
XFILLER_0_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10480__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net576 net577 vssd1 vssd1
+ vccd1 vccd1 _05652_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08339_ net2904 net2731 net1049 vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11350_ _07612_ _07613_ _05280_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__o21ai_1
X_10301_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] _04655_ vssd1
+ vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12543__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ net544 _07544_ _07542_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13020_ _06106_ _07807_ _07809_ _05549_ _07803_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__a221o_1
XANTENNA__09386__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10232_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\] net861 vssd1
+ vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__and3_1
XANTENNA__09925__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\] net859 vssd1
+ vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__and3_1
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10290__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1014 _04484_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__buf_2
Xfanout1025 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1025 sky130_fd_sc_hd__clkbuf_4
Xfanout1036 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1
+ net1036 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14131__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1052 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_14971_ net1298 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
X_10094_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] net888 vssd1
+ vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__and3_1
Xfanout1058 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1058 sky130_fd_sc_hd__clkbuf_2
Xfanout1069 net1071 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_1
X_16710_ clknet_leaf_129_wb_clk_i _02270_ _00573_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ net1167 net1059 net1790 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[3\]
+ sky130_fd_sc_hd__and3b_1
X_17690_ clknet_leaf_76_wb_clk_i _03250_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09153__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[27\]
+ _00504_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13853_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04113_ net1992 vssd1 vssd1
+ vccd1 vccd1 _04135_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10299__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14994__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ net3237 net199 net371 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16572_ clknet_leaf_142_wb_clk_i _02200_ _00435_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08992__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ _07707_ _04088_ net484 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__or3b_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10996_ _07164_ _07169_ net525 vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__mux2_2
XFILLER_0_35_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08113__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08113__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11799__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15523_ net1219 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12735_ net3058 net234 net379 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
XANTENNA__12718__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13403__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14198__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15454_ net1297 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
X_12666_ net2502 net209 net389 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14405_ net1308 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
X_11617_ net497 _07823_ net1948 net839 vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__o2bb2a_1
X_18173_ net1547 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
X_15385_ net1193 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
X_12597_ _07841_ _08012_ net488 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and3_4
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10465__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17124_ clknet_leaf_129_wb_clk_i _02684_ _00987_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11548_ _07705_ _07739_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__nand2_1
X_14336_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1 vssd1 vccd1
+ vccd1 _02262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold508 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold519 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[7\] vssd1 vssd1 vccd1 vccd1 net2135
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12453__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17055_ clknet_leaf_0_wb_clk_i _02615_ _00918_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] _04250_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\]
+ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ net319 _07701_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13218_ net2164 net2084 net818 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
X_16006_ net1358 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__inv_2
XANTENNA__09377__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\] _04275_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__a221o_1
XANTENNA__12920__A1 _07243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13149_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1208 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
X_17957_ clknet_leaf_106_wb_clk_i _03507_ _01777_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\]
+ sky130_fd_sc_hd__dfstp_1
Xhold1219 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
X_18176__1550 vssd1 vssd1 vccd1 vccd1 _18176__1550/HI net1550 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16908_ clknet_leaf_44_wb_clk_i _02468_ _00771_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11487__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17557__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ _04939_ _04940_ _04953_ net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__o32a_4
X_17888_ clknet_leaf_99_wb_clk_i _03438_ _01708_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16839_ clknet_leaf_121_wb_clk_i _02399_ _00702_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08104__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\] net705 _05572_
+ _05573_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12628__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14189__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\] net687 _05503_
+ _05504_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08407__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10656__B _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] net692 _05423_
+ _05427_ _05429_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_111_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout224_A _07915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ team_01_WB.instance_to_wrap.cpu.K0.code\[0\] _04552_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or3b_2
XFILLER_0_16_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10214__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09080__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08055_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 _04486_
+ sky130_fd_sc_hd__inv_2
XANTENNA__12363__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09907__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1300_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] net913
+ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__and3_1
XANTENNA__13194__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\] net704 _05139_
+ _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a211o_1
XANTENNA__08343__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10150__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09404__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _05515_ _05583_ net548 _05718_ net503 net518 vssd1 vssd1 vccd1 vccd1 _07114_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09701__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\] net727 _05763_ _05766_
+ _05770_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12538__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ _05166_ _05043_ net498 vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__mux2_1
XANTENNA__09843__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12520_ net2281 net262 net409 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__B2 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_137_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12451_ net2800 net246 net415 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ _07023_ _07665_ _07664_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10205__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15170_ net1290 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XANTENNA__11402__A1 _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ net2688 net280 net423 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13877__B team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09071__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14121_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\] _04278_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\]
+ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ _07054_ _07593_ _07595_ _07596_ _07591_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__a311o_1
XANTENNA__12273__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10582__A team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14052_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] _04149_ _04213_ vssd1
+ vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11264_ _06991_ _07073_ _07334_ _07061_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__o211a_1
XANTENNA__11166__B1 _07256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13003_ net2740 net217 net360 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10215_ _06475_ _06476_ _06477_ _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__or4_1
XANTENNA__16454__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11195_ _06384_ net343 vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__nand2_1
XANTENNA__08987__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17811_ clknet_leaf_68_wb_clk_i _03368_ _01632_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10146_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\] net734 _06392_ _06394_
+ _06399_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17742_ clknet_leaf_105_wb_clk_i _03300_ _01563_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10077_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\] net737 net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__a22o_1
X_14954_ net1201 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13905_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] net795 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[18\] sky130_fd_sc_hd__and2_1
X_17673_ clknet_leaf_73_wb_clk_i _03233_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14885_ net1312 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16624_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[10\]
+ _00487_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13836_ net1935 _04116_ _04127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[10\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13615__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16555_ clknet_leaf_93_wb_clk_i _02183_ _00418_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13767_ net1063 _07711_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__nor2_1
XANTENNA__13091__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12448__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10979_ _07226_ _07230_ _07242_ _07240_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__or4b_4
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ net1182 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
X_12718_ net2289 net263 net384 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XANTENNA__10444__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16486_ clknet_leaf_83_wb_clk_i _02114_ _00349_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_13698_ _04464_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18225_ net1588 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
X_15437_ net1216 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ net2673 net247 net391 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10195__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18156_ net1530 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
XANTENNA__13394__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ net1208 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XANTENNA__09984__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ clknet_leaf_48_wb_clk_i _02667_ _00970_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12183__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] _04455_ net1362 vssd1
+ vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold316 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ net1461 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_44_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15299_ net1209 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
Xhold327 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 _02009_ vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _01954_ vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09058__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17038_ clknet_leaf_53_wb_clk_i _02598_ _00901_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout807 _03743_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_8
X_09860_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] net954 vssd1
+ vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout818 net821 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_4
Xfanout829 net832 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
X_08811_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] _04657_
+ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and3_1
XANTENNA__16947__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\] net952 vssd1
+ vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__and3_1
Xhold1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] net633 net612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a22o_1
Xhold1038 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 team_01_WB.instance_to_wrap.cpu.f0.num\[20\] vssd1 vssd1 vccd1 vccd1 net2665
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] net639 net627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13082__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12358__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08628__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout439_A _08021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\] net948 vssd1
+ vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout606_A _03574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1348_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13385__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09156_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\] net962
+ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09894__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08107_ _04529_ _04533_ _04534_ _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__or4_1
XANTENNA__16477__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12093__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\] net949 vssd1
+ vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08038_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1 _04469_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold850 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 team_01_WB.instance_to_wrap.cpu.K0.code\[4\] vssd1 vssd1 vccd1 vccd1 net2477
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12821__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold883 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12896__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14602__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\] net732 net706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__a22o_1
XANTENNA__08564__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09761__B1 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08600__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] net963 vssd1
+ vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09513__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1550 _03454_ vssd1 vssd1 vccd1 vccd1 net3166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1561 _02049_ vssd1 vssd1 vccd1 vccd1 net3177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1572 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\] vssd1 vssd1 vccd1 vccd1
+ net3188 sky130_fd_sc_hd__dlygate4sd3_1
X_11951_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] net274 net472 vssd1
+ vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__mux2_1
XANTENNA__09134__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1583 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08867__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1594 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13652__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15433__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ net537 _07165_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11882_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__xor2_1
X_14670_ net1378 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09431__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ _07094_ _07096_ net526 vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__mux2_1
X_13621_ _07945_ _03956_ net188 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12268__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08619__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16340_ clknet_leaf_63_wb_clk_i net1858 _00208_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10426__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13552_ _03856_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10764_ net548 _05583_ net503 vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__mux2_1
XANTENNA__08047__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11623__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17252__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12503_ net2625 net202 net408 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
X_16271_ clknet_leaf_67_wb_clk_i _01908_ _00139_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ _03826_ _03828_ _03832_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ _06958_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18010_ clknet_leaf_79_wb_clk_i _03559_ _01824_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15222_ net1303 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
X_12434_ net3219 net190 net415 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13376__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15153_ net1199 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
X_12365_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] _07835_ _07840_ _07843_ vssd1
+ vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__and4b_1
XFILLER_0_80_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11316_ net545 _07560_ _07574_ _07080_ _07575_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__o221a_1
X_14104_ net792 _04237_ _04241_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__and3_4
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15084_ net1262 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12296_ net2028 net297 net434 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11139__A0 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14035_ net565 _04206_ _04207_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__and3_1
XANTENNA__15608__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ _05485_ _06037_ _06605_ _06870_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12731__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09606__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _06455_ _06594_ net345 vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08510__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] net932 vssd1
+ vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15986_ net1353 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__inv_2
XANTENNA__09504__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13300__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17725_ clknet_leaf_71_wb_clk_i _03283_ _01546_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14937_ net1237 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13562__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17656_ clknet_leaf_25_wb_clk_i _03216_ _01519_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14868_ net1339 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09341__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16607_ clknet_leaf_112_wb_clk_i _02235_ _00470_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08883__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ team_01_WB.instance_to_wrap.cpu.c0.count\[4\] team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17587_ clknet_leaf_49_wb_clk_i _03147_ _01450_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12178__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09807__B2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14799_ net1361 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16538_ clknet_leaf_59_wb_clk_i _02166_ _00401_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10417__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16469_ clknet_leaf_80_wb_clk_i _02097_ _00332_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11090__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09010_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\] net616 _05273_ net670
+ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17745__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ net1582 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
XANTENNA__13367__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09035__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ net1513 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 _01981_ vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold113 _03517_ vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold124 team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] vssd1 vssd1 vccd1 vccd1
+ net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold135 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 net1751
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold146 _01960_ vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 team_01_WB.instance_to_wrap.a1.ADR_I\[28\] vssd1 vssd1 vccd1 vccd1 net1773
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17895__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold168 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 net1784
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold179 net122 vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _06141_ _06175_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12641__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 net606 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_4
XFILLER_0_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12878__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout615 _04774_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_8
Xfanout626 _04766_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09843_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net591 net581 vssd1 vssd1
+ vccd1 vccd1 _06107_ sky130_fd_sc_hd__a21oi_1
Xfanout637 _04759_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_8
Xfanout648 net649 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08420__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _04739_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout389_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _05622_ _05761_ _06036_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__or3_1
XANTENNA__14095__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] net653 net622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1298_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11781__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\] net732 net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ _04908_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09889__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17275__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18235__1592 vssd1 vssd1 vccd1 vccd1 _18235__1592/HI net1592 sky130_fd_sc_hd__conb_1
XFILLER_0_117_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12088__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08587_ _04847_ _04850_ net580 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout723_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12816__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13358__A1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09208_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] net631 _05454_
+ _05461_ _05467_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a2111o_1
X_10480_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] net686 _06726_
+ _06729_ _06733_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__a2111o_1
X_18155__1529 vssd1 vssd1 vccd1 vccd1 _18155__1529/HI net1529 sky130_fd_sc_hd__conb_1
XFILLER_0_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09139_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\] net870
+ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12150_ net2821 net279 net448 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09129__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _06995_ _07352_ _07364_ net330 vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__a22o_1
X_12081_ net2774 net257 net456 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12551__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14332__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13530__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _05065_ net334 vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__nand2_1
XANTENNA__09426__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ net1287 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_139_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14086__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17618__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15771_ net1318 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ net1801 net604 net586 _03663_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17510_ clknet_leaf_137_wb_clk_i _03070_ _01373_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1380 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14722_ net1321 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1391 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3007 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11934_ net2832 net194 net473 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09161__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17441_ clknet_leaf_136_wb_clk_i _03001_ _01304_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14653_ net1369 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07849_ vssd1 vssd1 vccd1
+ vccd1 _07981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17768__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13597__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ _03829_ _03941_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_67_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10816_ net549 net543 net330 vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_32_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17372_ clknet_leaf_11_wb_clk_i _02932_ _01235_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14584_ net1396 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
X_11796_ net775 _07922_ _07923_ _07924_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__a2bb2o_4
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16323_ clknet_leaf_81_wb_clk_i net1702 _00191_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ net967 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] _03883_ _03884_
+ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a22o_1
XANTENNA__12726__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ _07007_ _07010_ net528 vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13349__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13411__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16254_ clknet_leaf_70_wb_clk_i _01891_ _00122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10678_ _06935_ _06941_ _04959_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__a21oi_1
X_13466_ _03817_ _03818_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16792__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15205_ net1232 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08225__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net2077 net276 net420 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
X_16185_ clknet_leaf_90_wb_clk_i _01853_ _00053_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13397_ net3194 net329 net353 team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1
+ vccd1 vccd1 _01886_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10473__C _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ net1273 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ net2541 net278 net491 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13539__A1_N net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17148__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net2449 net220 net431 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__mux2_1
X_15067_ net1315 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XANTENNA__12461__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14242__A _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09725__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\]
+ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__and3_2
XANTENNA__08878__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16172__CLK clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17298__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap890_A _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15969_ net1334 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__inv_2
XANTENNA__13285__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ net1077 net842 vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__and2_4
X_17708_ clknet_leaf_109_wb_clk_i _03268_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_09490_ _05720_ _05752_ net582 vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08441_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] net739 net734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ clknet_leaf_126_wb_clk_i _03199_ _01502_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09502__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08372_ _04624_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12636__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08415__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout304_A _07970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1046_A team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__C1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12371__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1213_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _03564_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_6
XANTENNA__09716__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 _03561_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_4
XANTENNA__08519__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16515__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13512__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 _08027_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_8
Xfanout434 _08023_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 _08020_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 net458 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout467 net470 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_8
X_09826_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] net893 vssd1
+ vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout478 _08009_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_6
Xfanout489 _08026_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_1
XANTENNA__13276__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\] net642 _04774_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\] vssd1 vssd1 vccd1 vccd1
+ _06021_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout840_A team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout938_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16665__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08708_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\] net752 net720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a22o_1
XANTENNA__11826__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ _05948_ _05949_ _05950_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__or4_1
XANTENNA__17910__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08639_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net763 net590 vssd1 vssd1
+ vccd1 vccd1 _04903_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ net1876 net1157 net567 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1
+ vccd1 vccd1 _03314_ sky130_fd_sc_hd__a22o_1
XANTENNA__09247__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14240__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ _06852_ _06861_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__nand2b_1
X_11581_ _07731_ _07794_ _07802_ net320 team_01_WB.instance_to_wrap.cpu.f0.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12546__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13320_ net134 net813 net807 net1723 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a22o_1
X_10532_ _06793_ _06794_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13251_ net59 net60 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__nand2_1
X_10463_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\] _04650_
+ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12202_ net3036 net190 net439 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XANTENNA_input67_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\] net636 net627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\]
+ _06647_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a221o_1
X_12133_ net3038 net210 net454 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
XANTENNA__08979__B net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12281__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ clknet_leaf_60_wb_clk_i _03539_ _01810_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16195__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12064_ net1865 net297 net462 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XANTENNA__09156__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16941_ clknet_leaf_21_wb_clk_i _02501_ _00804_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17440__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11514__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09183__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _07044_ _07048_ net510 vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16872_ clknet_leaf_61_wb_clk_i _02432_ _00735_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout990 net991 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_2
X_15823_ net1247 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13267__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13406__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15754_ net1198 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
X_12966_ net1033 _07414_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14705_ net1401 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ net2880 net217 net475 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
X_15685_ net1233 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
XANTENNA__09322__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11293__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12897_ net1620 net607 net589 _03601_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ clknet_leaf_25_wb_clk_i _02984_ _01287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10468__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ net1373 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
X_11848_ net2513 net264 net480 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14231__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ clknet_leaf_46_wb_clk_i _02915_ _01218_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08446__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ net1333 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12456__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ net775 _07908_ _07910_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__o21ai_4
XANTENNA__10253__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16306_ clknet_leaf_113_wb_clk_i _01940_ _00174_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ _07023_ _03870_ net767 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__mux2_1
X_17286_ clknet_leaf_141_wb_clk_i _02846_ _01149_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14498_ net1361 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16237_ clknet_leaf_79_wb_clk_i _00007_ _00105_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13449_ _03800_ _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16538__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16168_ clknet_leaf_57_wb_clk_i _01836_ _00036_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09992__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09410__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ net1248 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
XANTENNA__12191__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] net845
+ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__and3_1
X_16099_ net1400 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__inv_2
XANTENNA__09066__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08401__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16688__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17933__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[8\] net871 vssd1
+ vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18154__1528 vssd1 vssd1 vccd1 vccd1 _18154__1528/HI net1528 sky130_fd_sc_hd__conb_1
X_09542_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] net860 vssd1
+ vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09477__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__B _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08685__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\] net904 vssd1
+ vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__and3_1
XANTENNA__09232__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout254_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__B _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10492__B1 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ net1118 net940 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__and2_2
XFILLER_0_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14222__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08355_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] net1945 net1048 vssd1 vssd1
+ vccd1 vccd1 _03392_ sky130_fd_sc_hd__mux2_1
XANTENNA__11036__A2 _07185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08437__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1163_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10244__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ net2130 net2198 net1040 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1330_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13733__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout888_A _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1207 net1236 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_2
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout1218 net1236 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09407__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1229 net1235 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_4
Xfanout231 _07897_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_61_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout242 net245 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
Xfanout253 _07934_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout275 _07948_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_1
Xfanout286 net289 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
Xfanout297 _08001_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09704__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09809_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] net887 vssd1
+ vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ net1911 net243 net373 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12751_ net2866 net262 net382 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
XANTENNA__08676__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__D _07640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10288__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10483__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11702_ _07841_ _07842_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__nand2_1
X_15470_ net1230 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
X_12682_ net3000 net249 net388 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux2_1
X_14421_ net1282 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11633_ net1928 net840 _07808_ _07831_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__o22a_1
XANTENNA__13421__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12276__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17140_ clknet_leaf_6_wb_clk_i _02700_ _01003_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14352_ net1661 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11564_ _07701_ _07769_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nor2_1
XANTENNA__08055__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13303_ net121 net808 net803 net1877 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a22o_1
XANTENNA__17806__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13896__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10515_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\] net700 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a22o_1
X_17071_ clknet_leaf_18_wb_clk_i _02631_ _00934_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11495_ net483 _07725_ _07743_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__a21o_1
X_14283_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16022_ net1356 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__inv_2
X_10446_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] net655 _06709_
+ net670 vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__a211o_1
X_13234_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] net2227 net823 vssd1 vssd1
+ vccd1 vccd1 _02024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10377_ _06629_ _06634_ _06638_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13165_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
XANTENNA__08502__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12116_ net2134 net252 net452 vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__mux2_1
X_17973_ clknet_leaf_70_wb_clk_i _03522_ _01793_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13096_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\] net1028 vssd1 vssd1 vccd1
+ vccd1 _03718_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12047_ net2645 net221 net461 vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
XANTENNA__15616__A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16924_ clknet_leaf_15_wb_clk_i _02484_ _00787_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14520__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08903__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16980__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16855_ clknet_leaf_24_wb_clk_i _02415_ _00718_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15806_ net1315 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16786_ clknet_leaf_22_wb_clk_i _02346_ _00649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13998_ _04169_ _03553_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ net1193 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XANTENNA__09052__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\] _07510_ net1032 vssd1 vssd1
+ vccd1 vccd1 _03639_ sky130_fd_sc_hd__mux2_1
XANTENNA__08667__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10198__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10474__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15668_ net1241 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XANTENNA__09987__C _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14204__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17407_ clknet_leaf_1_wb_clk_i _02967_ _01270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14619_ net1363 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12186__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15599_ net1251 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08140_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04565_ vssd1 vssd1 vccd1 vccd1
+ _04567_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17338_ clknet_leaf_36_wb_clk_i _02898_ _01201_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17486__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08071_ net1748 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ sky130_fd_sc_hd__inv_2
X_17269_ clknet_leaf_8_wb_clk_i _02829_ _01132_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09919__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap965 _04638_ vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08412__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\] net735 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09227__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold17 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\] vssd1 vssd1 vccd1 vccd1 net1633
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold28 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\] vssd1 vssd1 vccd1 vccd1
+ net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A _04484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10701__A1 _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A _03571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] net667 vssd1 vssd1
+ vccd1 vccd1 _05789_ sky130_fd_sc_hd__nor2_2
XANTENNA__13651__A0 _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1280_A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A _04761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15261__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1378_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09456_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _05243_ _05242_ vssd1 vssd1
+ vccd1 vccd1 _05720_ sky130_fd_sc_hd__a21o_1
XANTENNA__09897__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16703__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ net1122 net921 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__and2_2
XANTENNA__12096__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] net762 _05649_ _05650_
+ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08338_ net2936 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ net2761 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[79\] net1045 vssd1 vssd1
+ vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
XANTENNA__12824__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08830__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] net939 vssd1
+ vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17979__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11280_ net538 _06991_ _07170_ _07335_ _07543_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__o311a_1
XFILLER_0_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] net843 vssd1
+ vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09386__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] net894 vssd1
+ vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 net1008 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09137__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1015 net1024 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13655__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1026 net1036 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_2
X_10093_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\] net883 vssd1
+ vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__and3_1
X_14970_ net1258 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
Xfanout1048 net1052 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14340__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09689__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1060 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_2
XANTENNA__12863__D_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09434__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ net1165 net1059 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[2\] sky130_fd_sc_hd__and3b_1
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16233__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17359__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[26\]
+ _00503_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ _04113_ _04134_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
X_12803_ net3230 net287 net371 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XANTENNA__12445__A1 _07925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16571_ clknet_leaf_5_wb_clk_i _02199_ _00434_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13783_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] _07706_ vssd1 vssd1 vccd1 vccd1
+ _04088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13642__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995_ _06955_ _07253_ _07258_ _06971_ _07257_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11903__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18225__1588 vssd1 vssd1 vccd1 vccd1 _18225__1588/HI net1588 sky130_fd_sc_hd__conb_1
XFILLER_0_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15522_ net1266 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
X_12734_ net2484 net202 net380 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18241_ net603 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
X_15453_ net1284 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
X_12665_ net2344 net193 net387 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
XANTENNA__09600__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14404_ net1308 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18172_ net1546 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
X_11616_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[18\] net573 vssd1 vssd1 vccd1
+ vccd1 _07823_ sky130_fd_sc_hd__nand2_1
X_15384_ net1254 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
X_12596_ net3253 net210 net402 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17123_ clknet_leaf_133_wb_clk_i _02683_ _00986_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14335_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1
+ vccd1 _02263_ sky130_fd_sc_hd__clkbuf_1
X_11547_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\] _07745_ _07778_ _07780_ vssd1
+ vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o211a_1
XANTENNA__12734__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10223__A3 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18153__1527 vssd1 vssd1 vccd1 vccd1 _18153__1527/HI net1527 sky130_fd_sc_hd__conb_1
XANTENNA__09609__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold509 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\] vssd1 vssd1 vccd1 vccd1
+ net2125 sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ clknet_leaf_4_wb_clk_i _02614_ _00917_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\] _04278_ _04280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\]
+ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11478_ net320 _07701_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__nor2_4
XANTENNA__08513__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16005_ net1355 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__inv_2
X_13217_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] net3176 net829 vssd1 vssd1
+ vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
X_10429_ _06690_ _06691_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11773__A1_N net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14197_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\] _04227_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\]
+ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13148_ net2993 net2607 net820 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XANTENNA__09047__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13565__S net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15346__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ net354 _03705_ _03706_ net834 net2382 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a32o_1
X_17956_ clknet_leaf_81_wb_clk_i net2353 _01776_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1209 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08886__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16907_ clknet_leaf_47_wb_clk_i _02467_ _00770_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_17887_ clknet_leaf_107_wb_clk_i net2509 _01707_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16838_ clknet_leaf_141_wb_clk_i _02398_ _00701_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ clknet_leaf_138_wb_clk_i _02329_ _00632_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\] net692 _05557_
+ _05561_ _05567_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10447__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\] net727 _05491_
+ _05493_ _05496_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a2111o_1
XANTENNA__16876__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08407__B net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\] net735 _05421_
+ _05426_ _05431_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08123_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\] team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11411__A2 _07669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout217_A _07943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10080__D1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08054_ net1120 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08423__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10672__B _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1126_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12911__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16256__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08956_ net978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] net947 vssd1
+ vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__and3_1
XANTENNA__17501__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] net703 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout753_A _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12427__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17651__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12819__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09508_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\] net915 vssd1
+ vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__and3_1
XANTENNA__10438__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _05241_ _05099_ net502 vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09439_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] net738 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11024__A _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12450_ net1973 net274 net416 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11401_ net1155 _04631_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12554__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12381_ net2438 net251 net425 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14335__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\] _04280_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a22o_1
X_11332_ net543 _06997_ _07173_ _07189_ _06955_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ _04213_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1
+ _04217_ sky130_fd_sc_hd__a31o_1
XANTENNA__11397__C _07659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ _05622_ net341 net337 _05621_ _07526_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11166__B2 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ net3133 net281 net362 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10214_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\] net693 _06460_ _06466_
+ _06468_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__a2111o_1
X_11194_ _06385_ _06595_ net345 vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__a21o_1
XANTENNA__13893__B net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\] _04651_ _04667_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] vssd1 vssd1 vccd1 vccd1
+ _06409_ sky130_fd_sc_hd__a22o_1
X_17810_ clknet_leaf_68_wb_clk_i _03367_ _01631_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17181__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09164__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16749__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17741_ clknet_leaf_96_wb_clk_i _03299_ _01562_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_14953_ net1205 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
X_10076_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\] net723 net717 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__a22o_1
X_13904_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] net795 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[17\] sky130_fd_sc_hd__and2_1
X_17672_ clknet_leaf_73_wb_clk_i _03232_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10103__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14884_ net1311 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
XANTENNA__10141__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16623_ clknet_leaf_96_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[9\]
+ _00486_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13835_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] _04116_ _04126_ vssd1 vssd1
+ vccd1 vccd1 _04127_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13414__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ clknet_leaf_55_wb_clk_i _02182_ _00417_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12969__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13766_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] _04014_ net1063 vssd1 vssd1 vccd1
+ vccd1 _04075_ sky130_fd_sc_hd__a21o_1
XANTENNA__13091__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10978_ net546 _07241_ _07079_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ net1192 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12717_ net2750 net266 net385 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
X_16485_ clknet_leaf_77_wb_clk_i _02113_ _00348_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09330__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] _04018_ vssd1 vssd1 vccd1 vccd1
+ _04019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18224_ net601 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
X_15436_ net1263 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
X_12648_ net2654 net277 net392 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13922__A_N net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18155_ net1529 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
XANTENNA__12464__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15367_ net1183 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
X_12579_ net2144 net250 net401 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__mux2_1
X_17106_ clknet_leaf_40_wb_clk_i _02666_ _00969_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14318_ _04455_ _04456_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18086_ net1460 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_124_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold306 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ net1286 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold317 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold328 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold339 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ clknet_leaf_18_wb_clk_i _02597_ _00900_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\] _04255_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[118\]
+ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11157__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_2
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout819 net820 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08573__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\] net914
+ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__and3_1
X_09790_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] net963 vssd1
+ vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__and3_1
XANTENNA__12106__A0 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] net628 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a22o_1
XANTENNA__17674__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17939_ clknet_leaf_83_wb_clk_i _03489_ _01759_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1028 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1039 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1390 net1398 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__buf_4
X_08672_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] net654 net613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12639__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09013__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11093__A0 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout334_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1076_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ _05349_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__or2_1
XANTENNA__09038__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17054__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12374__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _05378_ _05415_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08106_ _04462_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] team_01_WB.instance_to_wrap.cpu.f0.num\[22\]
+ _04467_ _04526_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09086_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] net963 vssd1
+ vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08037_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 _04468_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1410_A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold840 _02107_ vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold851 team_01_WB.instance_to_wrap.a1.ADR_I\[21\] vssd1 vssd1 vccd1 vccd1 net2467
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold873 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12896__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout870_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12896__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout968_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] net931 vssd1
+ vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10371__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08939_ _05166_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__and2_1
Xhold1540 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 net3156
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3167 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15714__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1562 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\] vssd1 vssd1 vccd1 vccd1
+ net3178 sky130_fd_sc_hd__dlygate4sd3_1
X_11950_ net2627 net217 net471 vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1573 _03448_ vssd1 vssd1 vccd1 vccd1 net3189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1584 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1595 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3211 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09712__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ _07161_ _07164_ net526 vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__mux2_1
X_18152__1526 vssd1 vssd1 vccd1 vccd1 _18152__1526/HI net1526 sky130_fd_sc_hd__conb_1
X_11881_ net3063 net311 net482 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__mux2_1
XANTENNA__12549__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ _03948_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ _07058_ _07095_ net516 vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13073__A1 _05549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13945__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14270__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11084__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ _03769_ _03852_ _03854_ _03855_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nand4_1
XFILLER_0_55_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10763_ _05923_ _05718_ net503 vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10831__A0 _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ net2678 net240 net408 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XANTENNA__09029__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16270_ clknet_leaf_68_wb_clk_i _01907_ _00138_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13482_ _03833_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__and2_1
X_10694_ _05043_ net498 _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15221_ net1173 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12433_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] _07869_ net417
+ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
XANTENNA__12284__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16421__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09159__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15152_ net1250 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12364_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] net213 net493 vssd1
+ vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14103_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\] _04263_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\]
+ _04262_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a221o_1
X_11315_ net321 _07578_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15083_ net1204 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
X_12295_ net2635 net308 net434 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14034_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\] _04147_ vssd1 vssd1 vccd1
+ vccd1 _04207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11246_ _07500_ _07501_ _07509_ _07499_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_30_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10898__A0 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13409__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11177_ _07430_ _07433_ _07440_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__and3b_2
XFILLER_0_78_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14089__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__B net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10128_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\] net939 vssd1
+ vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__and3_1
XANTENNA__09325__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15985_ net1381 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__inv_2
X_17724_ clknet_leaf_71_wb_clk_i _03282_ _01545_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10059_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\] net949 vssd1
+ vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__and3_1
X_14936_ net1254 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10114__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12459__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ net1339 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
X_17655_ clknet_leaf_12_wb_clk_i _03215_ _01518_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13818_ team_01_WB.instance_to_wrap.cpu.c0.count\[3\] team_01_WB.instance_to_wrap.cpu.c0.count\[2\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__and4_2
XFILLER_0_98_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ clknet_leaf_111_wb_clk_i _02234_ _00469_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_17586_ clknet_leaf_31_wb_clk_i _03146_ _01449_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14798_ net1308 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XANTENNA__14261__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17077__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16537_ clknet_leaf_62_wb_clk_i _02165_ _00400_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09060__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _07719_ _07774_ _04061_ net563 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10822__A0 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16468_ clknet_leaf_108_wb_clk_i _02096_ _00331_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09995__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15419_ net1299 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18207_ net1581 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
XANTENNA__12194__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16399_ clknet_leaf_75_wb_clk_i _02027_ _00262_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18138_ net1512 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
XFILLER_0_14_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16914__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold103 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\] vssd1 vssd1 vccd1 vccd1
+ net1719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10050__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold114 net114 vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold125 team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\] vssd1 vssd1 vccd1 vccd1
+ net1741 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ net1443 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__08794__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 _01970_ vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold147 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1 vccd1
+ net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold158 _02011_ vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ net582 _06174_ _06142_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__a21o_2
Xhold169 _01956_ vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12878__B2 _03587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout616 net617 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_8
X_09842_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__inv_2
Xfanout627 _04766_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout649 _04749_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_6
XANTENNA__10984__S0 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09773_ _05553_ _05621_ _06035_ _05552_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout284_A _07920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08724_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] net759 _04986_ _04987_
+ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09532__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] net752 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a22o_1
XANTENNA__12369__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout451_A _08018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1193_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net763 net590 vssd1 vssd1 vccd1
+ vccd1 _04850_ sky130_fd_sc_hd__a21o_1
XANTENNA__14252__B1 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout716_A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16444__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1360_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] net618 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13763__C1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\] net852
+ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16594__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08785__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] net903
+ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12832__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11100_ _04714_ _07211_ net531 vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09707__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ net2469 net220 net456 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
Xhold670 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold692 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13530__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ net532 _07072_ _07293_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13663__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ net1265 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _07441_ _03662_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] net1053
+ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1370 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08984__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ net1314 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11933_ _07841_ net495 _07846_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__and3_4
XANTENNA__12279__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1392 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] vssd1 vssd1 vccd1 vccd1
+ net3008 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17440_ clknet_leaf_141_wb_clk_i _03000_ _01303_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14652_ net1373 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
X_11864_ net2053 net242 net481 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14243__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13603_ _03826_ _03828_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__nand2_1
X_17371_ clknet_leaf_37_wb_clk_i _02931_ _01234_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13899__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10815_ _06990_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__and2_2
X_14583_ net1406 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\] net680 net775 vssd1 vssd1
+ vccd1 vccd1 _07924_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11911__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16322_ clknet_leaf_73_wb_clk_i net1785 _00190_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13534_ net771 _07640_ net967 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10746_ _07008_ _07009_ net518 vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16937__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16253_ clknet_leaf_71_wb_clk_i _01890_ _00121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13349__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _05653_ vssd1 vssd1
+ vccd1 vccd1 _03818_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10677_ _06934_ _06938_ _06940_ _06668_ _06939_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15204_ net1224 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ net2594 net217 net419 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__mux2_1
X_16184_ clknet_leaf_90_wb_clk_i _01852_ _00052_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ net2490 net328 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1
+ vccd1 vccd1 _01887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15135_ net1293 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
XANTENNA__08776__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ net2478 net251 net492 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11866__B _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15066_ net1257 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12278_ net2556 net283 net433 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__mux2_1
X_14017_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\] _04193_ vssd1 vssd1 vccd1
+ vccd1 _04194_ sky130_fd_sc_hd__and2_1
XANTENNA__08528__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ net534 net330 _07260_ _07333_ _07492_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__a311o_1
XFILLER_0_120_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08933__C1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09055__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11882__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15968_ net1336 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17707_ clknet_leaf_110_wb_clk_i _03267_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12189__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ net1184 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15899_ net1348 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08440_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\] net750 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ _04699_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a221o_1
X_17638_ clknet_leaf_136_wb_clk_i _03198_ _01501_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08371_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__nor3b_2
X_17569_ clknet_leaf_136_wb_clk_i _03129_ _01432_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08415__B _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12652__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18151__1525 vssd1 vssd1 vccd1 vccd1 _18151__1525/HI net1525 sky130_fd_sc_hd__conb_1
XFILLER_0_112_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09527__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08431__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10680__B _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 _03564_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_4
XANTENNA__08519__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 _03561_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 _08027_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout435 _08022_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout446 _08020_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17242__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_6
X_09825_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\] net865 vssd1
+ vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout479 net482 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_8
X_09756_ _06016_ _06017_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__or4_2
X_08707_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] net943
+ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__and3_1
XANTENNA__09262__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12099__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\] net640 _05926_ _05935_
+ _05941_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17392__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13028__A1 _03671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08638_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] net668 _04897_ _04901_
+ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o22a_4
XFILLER_0_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10201__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12827__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\] net656 net655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\]
+ _04830_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10600_ _06852_ _06863_ _06860_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__or3b_1
XFILLER_0_119_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11580_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] net1161 vssd1 vssd1 vccd1 vccd1
+ _07802_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10262__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10531_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\] net745 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__a22o_1
XANTENNA__10262__B2 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13250_ net56 net55 net58 net57 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10462_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] net918 vssd1
+ vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13658__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ net2235 net196 net441 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
XANTENNA__10014__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10014__B2 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10393_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] net625 _06656_ net672
+ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14343__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net2197 net292 net453 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__mux2_1
XANTENNA__09437__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16940_ clknet_leaf_48_wb_clk_i _02500_ _00803_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12063_ net1951 net307 net462 vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10317__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ _07276_ _07277_ net528 vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16871_ clknet_leaf_129_wb_clk_i _02431_ _00734_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11906__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 net993 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_2
X_15822_ net1217 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__inv_2
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08930__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15753_ net1215 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11278__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ net1623 net606 net588 _03650_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a22o_1
XANTENNA__11817__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ net1405 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
X_11916_ net2371 net279 net476 vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ net1272 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ net366 _03599_ _03600_ net1056 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ clknet_leaf_19_wb_clk_i _02983_ _01286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14635_ net1347 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XANTENNA__17885__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11847_ net778 _07964_ _07966_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12737__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14518__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13975__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ net1332 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
X_17354_ clknet_leaf_49_wb_clk_i _02914_ _01217_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ net681 _07307_ _07909_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16305_ clknet_leaf_113_wb_clk_i _01939_ _00173_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13517_ _07867_ _03869_ net186 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17285_ clknet_leaf_133_wb_clk_i _02845_ _01148_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ _04799_ net342 net333 _04798_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17115__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14497_ net1344 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16236_ clknet_leaf_34_wb_clk_i _00025_ _00104_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13448_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net592 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16167_ clknet_leaf_57_wb_clk_i _01835_ _00035_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12472__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ net2789 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1
+ vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10556__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15118_ net1234 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XANTENNA__12950__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17265__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16098_ net1388 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15049_ net1205 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_44_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\] net842 vssd1
+ vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__A _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\] net853 vssd1
+ vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10013__A1_N _06275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10021__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] net863 vssd1
+ vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14207__B1 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ net1118 net944 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__and2_2
XANTENNA__09810__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12647__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08354_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] net1939 net1048 vssd1 vssd1
+ vccd1 vccd1 _03393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08437__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08426__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08285_ net2939 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\] net1045 vssd1 vssd1
+ vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout414_A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11992__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17608__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13733__A2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12382__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10691__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1323_A net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10547__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09257__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16632__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 net212 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
Xfanout1208 net1211 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
Xfanout221 _07925_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout1219 net1227 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
Xfanout232 _07897_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
Xfanout243 net245 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net258 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
XANTENNA_fanout950_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 _07967_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout276 _07948_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout287 net289 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
X_09808_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] net858 vssd1
+ vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout298 net301 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16782__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] net881
+ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12750_ net1906 net267 net380 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09873__B1 _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11701_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12681_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] net274 net388 vssd1
+ vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XANTENNA__12557__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17138__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14338__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ net1280 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11632_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[10\] _07806_ vssd1 vssd1 vccd1
+ vccd1 _07831_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13421__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14351_ net3005 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__clkbuf_1
X_11563_ net320 _07788_ _07790_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13302_ net1795 net810 net805 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\] vssd1
+ vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a22o_1
XANTENNA__16162__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17070_ clknet_leaf_55_wb_clk_i _02630_ _00933_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10514_ _06776_ _06777_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__nor2_2
XANTENNA__17288__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14282_ net1778 _04201_ net1366 vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13896__B net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11494_ _07701_ _07740_ net319 vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_134_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16021_ net1355 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__inv_2
X_13233_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] net1720 net829 vssd1 vssd1
+ vccd1 vccd1 _02025_ sky130_fd_sc_hd__mux2_1
XANTENNA__12292__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\] net644 net635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__a22o_1
XANTENNA__11196__C1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09167__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13164_ net2869 net2718 net820 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10376_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\] net740 net690 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\]
+ _06639_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12115_ net3097 net256 net453 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17972_ clknet_leaf_70_wb_clk_i _03521_ _01792_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13095_ _05888_ _07807_ _03704_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__o21ai_1
X_16923_ clknet_leaf_38_wb_clk_i _02483_ _00786_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12046_ net1881 net285 net460 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13417__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16854_ clknet_leaf_29_wb_clk_i _02414_ _00717_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15805_ net1280 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09333__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13997_ _04181_ _04182_ _03556_ _04180_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__a2bb2o_1
X_16785_ clknet_leaf_23_wb_clk_i _02345_ _00648_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12948_ net2064 net605 net587 _03638_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15736_ net1257 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XANTENNA__09864__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18150__1524 vssd1 vssd1 vccd1 vccd1 _18150__1524/HI net1524 sky130_fd_sc_hd__conb_1
XANTENNA__09630__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11671__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ net1025 _07600_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__nand2_1
XANTENNA__12467__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15667_ net1187 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17406_ clknet_leaf_3_wb_clk_i _02966_ _01269_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14618_ net1410 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XANTENNA__09077__D1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15598_ net1228 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14549_ net1332 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17337_ clknet_leaf_16_wb_clk_i _02897_ _01200_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08070_ net1066 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17268_ clknet_leaf_7_wb_clk_i _02828_ _01131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16219_ clknet_leaf_42_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ _00087_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[0\] sky130_fd_sc_hd__dfrtp_1
Xmax_cap911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17199_ clknet_leaf_124_wb_clk_i _02759_ _01062_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10529__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17900__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11400__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09508__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14125__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\] net751 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__a22o_1
XANTENNA__10016__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09147__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 _02121_ vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14140__A2 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold29 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout197_A _07869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout364_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] net761 _05786_ _05787_
+ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__a22o_2
XANTENNA__15542__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09540__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] net576 net577 vssd1 vssd1
+ vccd1 vccd1 _05719_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12377__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1273_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout629_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ net1149 net1151 net1153 net1147 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__and4b_1
XANTENNA__16185__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] net710 net758 vssd1
+ vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17430__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11414__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08337_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] net1631 net1051 vssd1 vssd1
+ vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\] net2976 net1045 vssd1 vssd1
+ vccd1 vccd1 _03479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout998_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08199_ net1741 net553 _04568_ _04597_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17580__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13001__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10230_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\] net881 vssd1
+ vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09386__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__D1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10161_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\] net852 vssd1
+ vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__and3_1
XANTENNA__12840__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 net1008 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14131__A2 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1027 net1036 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
X_10092_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] net865 vssd1
+ vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__and3_1
Xfanout1038 net1046 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_2
Xfanout1049 net1052 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12142__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ net1166 net1059 net2370 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[1\]
+ sky130_fd_sc_hd__and3b_1
X_13851_ net2411 _04112_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nor2_1
XANTENNA__10299__C _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ net2720 net233 net373 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
X_13782_ net1693 _04087_ net782 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
X_16570_ clknet_leaf_3_wb_clk_i _02198_ _00433_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13642__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994_ _07177_ _07188_ net522 vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15521_ net1288 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
X_12733_ net2944 net240 net380 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
XANTENNA__12287__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11653__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18233__1591 vssd1 vssd1 vccd1 vccd1 _18233__1591/HI net1591 sky130_fd_sc_hd__conb_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15452_ net1279 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
X_18240_ net1593 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_12664_ net3255 _07869_ net389 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
XANTENNA__14198__A2 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14403_ net1351 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
X_11615_ net497 _07822_ net2190 net839 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__o2bb2a_1
X_18171_ net1545 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15383_ net1256 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12595_ net2500 net293 net402 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
XANTENNA__16678__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10759__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13700__A team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14334_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1
+ vccd1 _02264_ sky130_fd_sc_hd__clkbuf_1
X_17122_ clknet_leaf_143_wb_clk_i _02682_ _00985_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11546_ net1064 _07705_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1
+ vccd1 _07780_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ clknet_leaf_126_wb_clk_i _02613_ _00916_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\] _04227_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\]
+ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a22o_1
X_11477_ net483 _07729_ net320 vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16004_ net1406 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08513__B net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ net2329 net2178 net827 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\] net695 _06670_
+ _06671_ _06675_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09377__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14196_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\] _04233_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\]
+ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a22o_1
XANTENNA__09328__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15627__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ net2575 net1663 net824 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XANTENNA__12750__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10359_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\] net942
+ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__and3_1
XANTENNA__10392__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13078_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] net1028 vssd1 vssd1 vccd1
+ vccd1 _03706_ sky130_fd_sc_hd__or2_1
X_17955_ clknet_leaf_85_wb_clk_i net2284 _01775_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12029_ net2535 net311 net465 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
X_16906_ clknet_leaf_48_wb_clk_i _02466_ _00769_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17303__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17886_ clknet_leaf_98_wb_clk_i _03436_ _01706_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16837_ clknet_leaf_131_wb_clk_i _02397_ _00700_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09063__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16768_ clknet_leaf_141_wb_clk_i _02328_ _00631_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17453__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09360__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15719_ net1184 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XANTENNA__12197__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16699_ clknet_leaf_30_wb_clk_i _02259_ _00562_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09240_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\] net695 _05489_
+ _05498_ net711 vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14189__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09171_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] net689 _05420_
+ _05425_ _05430_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_84_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08122_ team_01_WB.instance_to_wrap.cpu.K0.code\[6\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__or4b_2
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08704__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ net1086 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11250__A1_N net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08423__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08576__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1021_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10383__B1 _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09535__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] net941
+ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08886_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\] net945
+ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1390_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13624__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] net739 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a22o_1
XANTENNA__09270__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09701__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17946__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09438_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] net940 vssd1
+ vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] net953
+ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__and3_1
XANTENNA__12835__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _04631_ vssd1 vssd1 vccd1
+ vccd1 _07664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ net2041 net256 net423 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16970__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ net527 _07594_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14050_ net2889 _04215_ _04216_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11262_ _05583_ _05620_ net331 _07525_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_127_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11166__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08567__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ net2605 net252 net361 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
X_10213_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\] net727 _06458_ _06464_
+ _06467_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13666__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12570__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _06385_ _06879_ _06884_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__nor3_1
XANTENNA_input42_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08987__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _06397_ _06405_ _06406_ _06407_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11186__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17740_ clknet_leaf_104_wb_clk_i net1870 _01561_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10075_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] net754 _06322_ _06323_
+ _06327_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__a2111o_1
X_14952_ net1181 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] net795 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[16\] sky130_fd_sc_hd__and2_1
X_17671_ clknet_leaf_123_wb_clk_i _03231_ _01534_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14883_ net1311 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11914__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16622_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[8\]
+ _00485_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13834_ _04120_ _04121_ _04126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13615__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13765_ net1654 net782 _04073_ _04074_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16553_ clknet_leaf_20_wb_clk_i _02181_ _00416_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10977_ net539 _07134_ _07234_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09611__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15504_ net1256 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12716_ net1946 net270 net383 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13696_ net1062 _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__or2_1
X_16484_ clknet_leaf_108_wb_clk_i _02112_ _00347_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18223_ net602 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15435_ net1210 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
X_12647_ net2389 net217 net391 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XANTENNA__12745__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11929__A1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13430__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18154_ net1528 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
X_15366_ net1287 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12578_ net3066 net254 net399 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ clknet_leaf_24_wb_clk_i _02665_ _00968_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11529_ net483 _07765_ net319 vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__a21o_1
X_14317_ net1884 _04454_ net1172 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__o21ai_1
X_15297_ net1312 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
X_18085_ net1459 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
Xhold307 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\] vssd1 vssd1 vccd1 vccd1
+ net1934 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ clknet_leaf_47_wb_clk_i _02596_ _00899_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold329 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[1\] vssd1 vssd1 vccd1 vccd1
+ net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] _04227_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\]
+ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09058__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15357__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14179_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\] _04272_ _04275_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\]
+ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__a221o_1
XANTENNA__12480__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net811 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
X_08740_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] net642 net629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a22o_1
X_17938_ clknet_leaf_78_wb_clk_i net2802 _01758_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1018 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\] vssd1 vssd1 vccd1 vccd1
+ net2634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10668__A1 _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1380 net1389 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__buf_4
Xfanout1391 net1398 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__buf_2
X_08671_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] net759 _04933_ _04934_
+ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a22o_2
X_17869_ clknet_leaf_104_wb_clk_i _03419_ _01689_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08730__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15092__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17969__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10948__B _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09286__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11093__A1 _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ _05419_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12655__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1069_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ _05378_ _05416_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nor2_1
X_08105_ _04461_ team_01_WB.instance_to_wrap.cpu.f0.num\[30\] team_01_WB.instance_to_wrap.cpu.f0.num\[25\]
+ _04464_ _04513_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_115_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08797__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16223__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13790__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09085_ _05281_ _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1236_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08036_ team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1 _04467_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold830 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold841 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold852 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12390__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 team_01_WB.instance_to_wrap.cpu.f0.num\[2\] vssd1 vssd1 vccd1 vccd1 net2490
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1403_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\] vssd1 vssd1 vccd1 vccd1
+ net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09265__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17499__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] _04657_
+ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout863_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08600__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net578 _05199_ _05200_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__o21a_1
XANTENNA__10204__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1530 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09513__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1541 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3168 sky130_fd_sc_hd__dlygate4sd3_1
X_08869_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] net666 _05127_ _05132_
+ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__o22a_4
XFILLER_0_58_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16098__A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1563 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1574 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 net3190
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1585 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3201 sky130_fd_sc_hd__dlygate4sd3_1
X_10900_ _07162_ _07163_ net514 vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__mux2_1
XANTENNA__08721__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1596 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\] vssd1 vssd1 vccd1 vccd1
+ net3212 sky130_fd_sc_hd__dlygate4sd3_1
X_11880_ _07992_ _07993_ net778 vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__mux2_4
XFILLER_0_93_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10831_ _04883_ _04935_ net498 vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09431__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _03895_ _03896_ net1066 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10762_ net322 _07025_ _06947_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ net1988 net208 net407 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10831__A1 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _05310_ vssd1 vssd1
+ vccd1 vccd1 _03834_ sky130_fd_sc_hd__xor2_1
X_10693_ _04988_ net498 vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12565__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14346__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15220_ net1242 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
X_12432_ _07846_ _08008_ net488 vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11387__A2 _07258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15151_ net1248 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
X_12363_ net2578 net293 net491 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
X_14102_ net788 _04237_ _04241_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__and3_4
X_11314_ _07576_ _07577_ net533 vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15082_ net1197 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
X_12294_ net2274 net312 net434 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14033_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\] _04147_ vssd1 vssd1 vccd1
+ vccd1 _04206_ sky130_fd_sc_hd__or2_1
XANTENNA__11909__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ net547 _07508_ _07507_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09752__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ net547 _07427_ _07439_ _07107_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09606__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] _04655_
+ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__and3_1
XANTENNA__15905__A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15984_ net1381 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17723_ clknet_leaf_71_wb_clk_i team_01_WB.instance_to_wrap.cpu.K0.next_keyvalid
+ _01544_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.keyvalid sky130_fd_sc_hd__dfrtp_4
XANTENNA__09504__A2 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] net946 vssd1
+ vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14935_ net1238 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08712__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17654_ clknet_leaf_30_wb_clk_i _03214_ _01517_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14866_ net1339 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16605_ clknet_leaf_118_wb_clk_i _02233_ _00468_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13817_ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__nand2_1
XANTENNA__09341__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17585_ clknet_leaf_20_wb_clk_i _03145_ _01448_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14797_ net1394 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_69_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16536_ clknet_leaf_64_wb_clk_i _02164_ _00399_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13748_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] team_01_WB.instance_to_wrap.cpu.f0.i\[19\]
+ _04015_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 _04061_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10822__A1 _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16467_ clknet_leaf_100_wb_clk_i _02095_ _00330_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_13679_ net772 _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18206_ net1580 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
XFILLER_0_5_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15418_ net1265 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ clknet_leaf_82_wb_clk_i _02026_ _00261_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08779__B1 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18137_ net1511 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
XANTENNA__13772__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15349_ net1173 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold104 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\] vssd1 vssd1 vccd1 vccd1 net1720
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold115 _01966_ vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10050__A2 _06313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16396__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold126 team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\] vssd1 vssd1 vccd1 vccd1
+ net1742 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ net1442 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17641__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold137 net99 vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold148 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\] vssd1 vssd1 vccd1 vccd1
+ net1764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11819__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold159 team_01_WB.instance_to_wrap.a1.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 net1775
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ clknet_leaf_32_wb_clk_i _02579_ _00882_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09910_ _06169_ _06171_ _06173_ _06143_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__o31a_2
XFILLER_0_121_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12878__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 _03574_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_4
Xfanout617 _04773_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_8
XFILLER_0_95_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] net667 _06101_ _06104_
+ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__o22ai_4
XANTENNA__10889__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 _04765_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_8
Xfanout639 _04758_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_8
XANTENNA__08420__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _05515_ _05551_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__xnor2_4
XANTENNA__17791__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] net698 net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10510__A0 _06772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08429__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17021__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08585_ net781 net765 _04715_ net682 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o41a_1
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout444_A _08020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1186_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12385__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout611_A _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17171__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09206_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\] net638 net633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\]
+ _05462_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a221o_1
XANTENNA__16739__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09137_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] net879
+ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10041__A2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[18\] net851 vssd1
+ vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout980_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11729__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1 vccd1 net2298
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net531 _07060_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__o21ai_1
Xhold693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09426__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ net1027 net364 vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] vssd1 vssd1 vccd1 vccd1
+ net2976 sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ net1320 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1371 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2987 sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ net2991 net212 net478 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__mux2_1
Xhold1382 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 _02134_ vssd1 vssd1 vccd1 vccd1 net3009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11863_ net778 _07977_ _07978_ _07979_ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__a2bb2o_1
X_14651_ net1347 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XANTENNA__16269__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17514__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13602_ net966 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _03939_ _03940_
+ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
X_10814_ net546 _06992_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__nand2_1
X_17370_ clknet_leaf_35_wb_clk_i _02930_ _01233_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14582_ net1347 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
X_11794_ net676 _07625_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__nand2_1
XANTENNA__13899__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16321_ clknet_leaf_73_wb_clk_i net1724 _00189_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12295__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13533_ net771 _03882_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__or2_1
X_10745_ _05993_ _05923_ net504 vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16252_ clknet_leaf_79_wb_clk_i _01889_ _00120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13464_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] _05653_ vssd1 vssd1
+ vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand2_1
X_10676_ _06718_ _06697_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17664__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15203_ net1220 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
X_12415_ net2345 net278 net420 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13395_ net3203 net327 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1
+ vccd1 vccd1 _01888_ sky130_fd_sc_hd__a22o_1
X_16183_ clknet_leaf_90_wb_clk_i _01851_ _00051_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09422__A1 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12346_ net2013 net256 net490 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__mux2_1
X_15134_ net1300 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09973__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__A _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11639__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15065_ net1190 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_116_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12277_ net2322 net222 net433 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__mux2_1
X_14016_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _04193_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09725__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _06997_ _07251_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__and2_1
XANTENNA__09336__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11159_ _06856_ _06867_ _06888_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__and3_1
XANTENNA__12978__B net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11882__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15967_ net1334 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__inv_2
XANTENNA__09489__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13285__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17706_ clknet_leaf_110_wb_clk_i _03266_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14918_ net1271 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15898_ net1348 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08161__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17637_ clknet_leaf_135_wb_clk_i _03197_ _01500_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14849_ net1353 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XANTENNA__17194__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _04624_ _04633_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__and2_1
X_17568_ clknet_leaf_141_wb_clk_i _03128_ _01431_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12796__A1 _07869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11143__S1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16519_ clknet_leaf_75_wb_clk_i _02147_ _00382_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17499_ clknet_leaf_37_wb_clk_i _03059_ _01362_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10559__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14714__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11756__C1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08431__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09177__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14170__B1 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13935__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 _03563_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_6
Xfanout414 _03561_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout425 _08027_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_6
XANTENNA_fanout394_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 _08022_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_4
XANTENNA__08924__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout447 _08019_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_6
X_09824_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] net848 vssd1
+ vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1101_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 _08016_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_6
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09543__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\] net663 _06006_
+ _06008_ _06012_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout659_A _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] net929
+ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__and3_1
XANTENNA__11287__A1 _06869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\] net643 _05928_
+ _05938_ _05946_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08152__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08637_ _04886_ _04887_ _04899_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or4_1
XFILLER_0_136_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout826_A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08568_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] net650 net624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\]
+ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16561__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08499_ net1084 net861 vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__and2_2
XFILLER_0_119_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13004__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10530_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\] net742 _06785_
+ _06788_ _06789_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_9_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11032__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] net913 vssd1
+ vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12843__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12200_ _07841_ net494 _08017_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ net2812 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] net820 vssd1 vssd1
+ vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XANTENNA__11967__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10392_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] net643 net637 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12131_ net3043 net296 net454 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09168__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17067__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net2817 net311 net462 vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XANTENNA__14161__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold490 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09156__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12711__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _07030_ _07035_ net512 vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16870_ clknet_leaf_141_wb_clk_i _02430_ _00733_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10183__D1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10722__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08995__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15821_ net1212 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__inv_2
Xfanout981 net993 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13267__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15752_ net1197 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
X_12964_ net365 _03648_ _03649_ net1055 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08143__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_115_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14703_ net1372 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ net2201 net251 net477 vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ net1223 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
X_12895_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1
+ vccd1 _03600_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11922__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17422_ clknet_leaf_53_wb_clk_i _02982_ _01285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ net1401 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ net681 _07510_ _07965_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11125__S1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ clknet_leaf_39_wb_clk_i _02913_ _01216_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14565_ net1331 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08446__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11777_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\] net674 net777 vssd1 vssd1
+ vccd1 vccd1 _07909_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11416__A2_N _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16304_ clknet_leaf_115_wb_clk_i _01938_ _00172_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10253__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13516_ _03867_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__xnor2_1
X_10728_ _04714_ net330 vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17284_ clknet_leaf_128_wb_clk_i _02844_ _01147_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14496_ net1362 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ clknet_leaf_42_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\]
+ _00103_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12753__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13447_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ net592 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__nand3_1
X_10659_ _05277_ _05241_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10005__A2 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13378_ net2665 net328 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1
+ vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
X_16166_ clknet_leaf_57_wb_clk_i _01834_ _00034_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12950__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15117_ net1216 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
X_12329_ net1995 net294 net430 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16097_ net1372 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14152__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15048_ net1204 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XANTENNA__09066__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16434__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10713__B1 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09363__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16999_ clknet_leaf_126_wb_clk_i _02559_ _00862_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] net848 vssd1
+ vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10302__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11117__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\] net896
+ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08685__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] net952 vssd1
+ vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10492__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__D1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08707__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] net1649 net1048 vssd1 vssd1
+ vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08437__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08426__B _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08284_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] net2401 net1041 vssd1 vssd1
+ vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1051_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09538__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_70_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10691__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10952__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1316_A net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14143__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_1
XFILLER_0_121_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1209 net1211 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
Xfanout233 _07897_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_1
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xfanout255 net258 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout266 net269 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_2
XANTENNA__09273__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 _07948_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
X_09807_ net555 _06070_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] net762
+ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__a2bb2o_4
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
XANTENNA__09704__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 net301 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout943_A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09738_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\] net867
+ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09669_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\] net866
+ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__and3_1
XANTENNA__08676__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11700_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__nor2_2
XANTENNA__10483__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12680_ net2238 net215 net387 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08617__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ net1952 net840 _07808_ _07830_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11562_ _07723_ _07734_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1
+ vccd1 _07790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11432__A1 _04593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14350_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1 vssd1 vccd1
+ vccd1 _02248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13301_ net1857 net808 net803 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\] vssd1
+ vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10513_ _06752_ _06774_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14281_ net1639 net1170 _04158_ _04434_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a31o_1
X_11493_ _07725_ _07741_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12573__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16020_ net1410 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__inv_2
X_13232_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] net2279 net827 vssd1 vssd1
+ vccd1 vccd1 _02026_ sky130_fd_sc_hd__mux2_1
XANTENNA_input72_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\] net648 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\]
+ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11196__B1 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12932__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ net2715 net2685 net824 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10375_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] net736 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10943__A0 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ net3024 net221 net453 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__mux2_1
XANTENNA__14134__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13094_ net354 _03715_ _03716_ net835 net2786 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a32o_1
X_17971_ clknet_leaf_78_wb_clk_i _03520_ _01791_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.InstrRead
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11917__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16922_ clknet_leaf_36_wb_clk_i _02482_ _00785_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12045_ net2293 net225 net459 vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
XANTENNA__09010__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18099__1473 vssd1 vssd1 vccd1 vccd1 _18099__1473/HI net1473 sky130_fd_sc_hd__conb_1
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13417__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16853_ clknet_leaf_26_wb_clk_i _02413_ _00716_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15804_ net1234 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16784_ clknet_leaf_25_wb_clk_i _02344_ _00647_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08116__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13996_ net1170 _04159_ _04163_ _03556_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a31o_1
XANTENNA__09313__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ net1238 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
X_12947_ net364 _03636_ _03637_ net1054 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__a32o_1
XANTENNA__12748__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08667__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10474__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15666_ net1178 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
X_12878_ net1836 net607 net589 _03587_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a22o_1
XANTENNA__11671__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17405_ clknet_leaf_14_wb_clk_i _02965_ _01268_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14617_ net1400 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11829_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\] _07551_ net679 vssd1 vssd1
+ vccd1 vccd1 _07952_ sky130_fd_sc_hd__mux2_1
X_15597_ net1218 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17336_ clknet_leaf_29_wb_clk_i _02896_ _01199_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14548_ net1331 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17232__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17267_ clknet_leaf_50_wb_clk_i _02827_ _01130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_131_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14479_ net1393 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16218_ clknet_leaf_71_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_atmax _00086_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.enable sky130_fd_sc_hd__dfrtp_1
XANTENNA__09358__A _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09919__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap901 net902 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_2
X_17198_ clknet_leaf_52_wb_clk_i _02758_ _01061_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12923__A1 _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap934 _04663_ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16149_ net1322 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__inv_2
XANTENNA__17382__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14125__B1 _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08971_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] net727 _05232_
+ _05233_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold19 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[10\] vssd1 vssd1 vccd1 vccd1
+ net1635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09552__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10032__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13100__A1 _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09304__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] net709 net757 vssd1
+ vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09821__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12658__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout357_A _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] net759 _05716_ _05717_
+ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__a22o_4
XANTENNA_fanout1099_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08405_ net971 net924 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ _05638_ _05640_ _05645_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__or4_4
XFILLER_0_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1266_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10217__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08336_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08871__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11798__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ net3128 net3094 net1049 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
XANTENNA__12393__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08830__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09268__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _04566_ _04596_ vssd1 vssd1 vccd1
+ vccd1 _04597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11178__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14902__A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\] net859 vssd1
+ vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17875__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1017 net1024 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_2
X_10091_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] net908 vssd1
+ vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__and3_1
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1039 net1041 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09434__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08897__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15733__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850_ _04112_ _04126_ _04133_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[5\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_134_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09731__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ net2951 net235 net371 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13781_ net484 _07709_ _07768_ _04086_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__a31o_1
XANTENNA__12568__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ _05418_ _07255_ _07256_ _07185_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__a2bb2o_1
X_15520_ net1286 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
XANTENNA__14009__A_N net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ net2540 net209 net380 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11653__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17255__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10596__B net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15451_ net1317 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12663_ _07845_ _08017_ net489 vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and3_4
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14402_ net1351 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
X_18170_ net1544 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
X_11614_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[19\] net573 vssd1 vssd1 vccd1
+ vccd1 _07822_ sky130_fd_sc_hd__nand2_1
X_15382_ net1303 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12594_ net2321 net295 net402 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XANTENNA__09074__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17121_ clknet_leaf_136_wb_clk_i _02681_ _00984_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14333_ net3033 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] _07778_ _07779_ _07731_ vssd1
+ vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08821__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17052_ clknet_leaf_15_wb_clk_i _02612_ _00915_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11476_ _04462_ _04505_ _07703_ _07727_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__or4b_1
X_14264_ _04414_ _04416_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or3_1
XANTENNA__08082__A _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09609__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16003_ net1386 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__inv_2
XANTENNA__12905__A1 _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13215_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\] net2431 net830 vssd1 vssd1
+ vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
X_10427_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] net697 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14195_ net1171 _04352_ _04353_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__and3_1
XANTENNA__08585__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\] net921
+ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__and3_1
X_13146_ net2636 net2571 net820 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
XANTENNA__08810__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10392__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13428__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17954_ clknet_leaf_79_wb_clk_i _03504_ _01774_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_13077_ net559 _07807_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__o21ai_1
X_10289_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] net621 _06550_ _06551_
+ _06552_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16905_ clknet_leaf_40_wb_clk_i _02465_ _00768_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12028_ net2093 net261 net466 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11341__A0 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17885_ clknet_leaf_104_wb_clk_i _03435_ _01705_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_79_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08888__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16836_ clknet_leaf_129_wb_clk_i _02396_ _00699_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09641__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12478__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13094__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ clknet_leaf_5_wb_clk_i _02327_ _00630_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13979_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[4\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ net584 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15718_ net1274 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10447__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ clknet_leaf_31_wb_clk_i _02258_ _00561_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ net1288 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16622__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09170_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] net695 _05422_
+ _05424_ _05428_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08121_ _04540_ _04542_ _04544_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ clknet_leaf_130_wb_clk_i _02879_ _01182_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13102__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] vssd1 vssd1 vccd1 vccd1
+ _04483_ sky130_fd_sc_hd__inv_2
XANTENNA__09088__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17898__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16772__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10027__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09816__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08954_ net978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\] net928 vssd1
+ vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1014_A _04484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08885_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\] net925 vssd1
+ vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__and3_1
XANTENNA__09254__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A _08010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15553__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10540__D1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17278__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1383_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\] net955 vssd1
+ vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__and3_1
XANTENNA__10438__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ net973 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] net929 vssd1
+ vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13801__A team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13388__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09368_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] net935
+ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__and3_1
X_18098__1472 vssd1 vssd1 vccd1 vccd1 _18098__1472/HI net1472 sky130_fd_sc_hd__conb_1
XFILLER_0_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08319_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09299_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] net943
+ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13012__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10071__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11330_ _06965_ _06975_ net510 vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11261_ _05620_ net335 vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__nand2_1
XANTENNA__15728__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12851__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12899__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13000_ net2956 net256 net362 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
X_10212_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\] net730 _04685_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a22o_1
XANTENNA__13560__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _07448_ _07455_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13248__A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\] net716 net694 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\] net722 _06320_ _06325_
+ _06330_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__a2111o_1
X_14951_ net1184 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XANTENNA__09164__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13902_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] net797 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[15\] sky130_fd_sc_hd__and2_1
X_17670_ clknet_leaf_139_wb_clk_i _03230_ _01533_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ net1311 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XANTENNA__10103__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ clknet_leaf_98_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[7\]
+ _00484_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13833_ team_01_WB.instance_to_wrap.cpu.c0.count\[16\] _04111_ _04124_ _04125_ vssd1
+ vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__nand4_2
XFILLER_0_76_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12298__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16552_ clknet_leaf_45_wb_clk_i _02180_ _00415_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ net484 _07715_ _07760_ net786 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__a31o_1
X_10976_ _07139_ _07186_ _07239_ net546 _07236_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15503_ net1202 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XANTENNA__11215__B _07441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12715_ net1897 net247 net384 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
X_16483_ clknet_leaf_100_wb_clk_i _02111_ _00346_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13695_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] _07718_ _07773_ team_01_WB.instance_to_wrap.cpu.f0.i\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11930__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18222_ net601 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13379__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15434_ net1197 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
X_12646_ net2922 net281 net392 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16795__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08805__A _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18153_ net1527 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
XANTENNA__13430__B _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15365_ net1222 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12577_ net3238 net220 net399 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17104_ clknet_leaf_25_wb_clk_i _02664_ _00967_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\] _04454_ vssd1 vssd1 vccd1
+ vccd1 _04455_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ _07708_ _07739_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__nand2_1
X_18084_ net1458 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
X_15296_ net1276 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09339__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold308 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 team_01_WB.instance_to_wrap.cpu.c0.count\[10\] vssd1 vssd1 vccd1 vccd1 net1935
+ sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ clknet_leaf_46_wb_clk_i _02595_ _00898_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12761__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\] _04239_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\]
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a22o_1
X_11459_ _07711_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__inv_2
XANTENNA__18014__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09636__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\] _04229_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\]
+ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08540__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13129_ net2542 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\] net828 vssd1 vssd1
+ vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16175__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09507__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ clknet_leaf_101_wb_clk_i _03487_ _01757_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15373__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1370 net1414 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__clkbuf_2
X_08670_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__o21a_1
X_17868_ clknet_leaf_75_wb_clk_i net1918 _01688_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1381 net1389 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__clkbuf_4
Xfanout1392 net1398 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16819_ clknet_leaf_49_wb_clk_i _02379_ _00682_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_17799_ clknet_leaf_59_wb_clk_i _03356_ _01620_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10310__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11617__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14717__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09038__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09153_ _05378_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] _04490_ team_01_WB.instance_to_wrap.cpu.f0.num\[23\]
+ _04466_ _04527_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _05346_ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ net1062 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15548__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold820 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12671__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1131_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold831 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold842 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold853 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16518__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold864 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\] vssd1 vssd1 vccd1 vccd1
+ net2480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09210__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold886 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12896__A3 _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold897 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09986_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] net932 vssd1
+ vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08937_ net578 _05199_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_23_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout856_A _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1520 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3158 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11856__A1 _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1553 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17913__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _05128_ _05129_ _05130_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or4_1
Xhold1564 team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\] vssd1 vssd1 vccd1 vccd1
+ net3180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1575 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1586 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 net3202
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09712__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1597 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[25\] vssd1 vssd1 vccd1 vccd1
+ net3213 sky130_fd_sc_hd__dlygate4sd3_1
X_08799_ net562 net561 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] net666
+ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__o2bb2a_4
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13007__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10830_ _07092_ _07093_ net514 vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09277__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14270__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12846__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ _04854_ _06943_ _06946_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ net3016 net192 net407 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09029__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10692_ _05099_ _05166_ net500 vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__mux2_1
X_13480_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] _05244_ vssd1 vssd1
+ vccd1 vccd1 _03833_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12033__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ net2934 net213 net422 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
XANTENNA__13230__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15150_ net1216 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ net2610 net294 net493 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09159__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11792__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101_ net792 net791 _04232_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__and3_4
X_11313_ _06960_ _06976_ net520 vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15081_ net1212 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
XANTENNA__12581__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12293_ net1896 net259 net433 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14032_ _04148_ net565 _04205_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__and3_1
XANTENNA__08998__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11244_ net330 _07135_ _07142_ _07333_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net541 _07438_ _07437_ _07436_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14089__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] net959 vssd1
+ vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ net1385 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__inv_2
X_17722_ clknet_leaf_71_wb_clk_i team_01_WB.instance_to_wrap.cpu.K0.next_state _01543_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.state sky130_fd_sc_hd__dfrtp_1
XANTENNA__11925__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] net949 vssd1
+ vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__and3_1
XANTENNA__13706__A team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11847__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14934_ net1259 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ clknet_leaf_25_wb_clk_i _03213_ _01516_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14865_ net1339 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16604_ clknet_leaf_112_wb_clk_i _02232_ _00467_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13816_ net2115 net785 _04559_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1
+ vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
XANTENNA__10130__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17584_ clknet_leaf_25_wb_clk_i _03144_ _01447_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14796_ net1354 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14261__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16535_ clknet_leaf_62_wb_clk_i _02163_ _00398_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13747_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] _07718_ vssd1 vssd1 vccd1 vccd1
+ _04060_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10959_ net324 _07219_ _07222_ _07218_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__o211a_2
XFILLER_0_112_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13441__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16466_ clknet_leaf_108_wb_clk_i _02094_ _00329_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13678_ _07995_ _04002_ net187 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18205_ net1579 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
XFILLER_0_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15417_ net1192 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ net2952 net212 net398 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XANTENNA__08228__B1 _00020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16397_ clknet_leaf_73_wb_clk_i _02025_ _00260_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08779__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18136_ net1510 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_38_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15348_ net1240 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09069__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09440__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11783__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18067_ net1441 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold105 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\] vssd1 vssd1 vccd1 vccd1
+ net1721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\] vssd1 vssd1 vccd1 vccd1
+ net1732 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ net1249 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[31\] vssd1 vssd1 vccd1 vccd1
+ net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold138 _02014_ vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ clknet_leaf_34_wb_clk_i _02578_ _00881_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13524__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09366__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\] vssd1 vssd1 vccd1 vccd1
+ net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09840_ _06095_ _06096_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__or4_2
Xfanout607 _03574_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 _04771_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10305__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17936__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13288__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ _05622_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__or2_1
X_18097__1471 vssd1 vssd1 vccd1 vccd1 _18097__1471/HI net1471 sky130_fd_sc_hd__conb_1
X_08722_ _04977_ _04979_ _04983_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__or4_4
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16960__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\] net938
+ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__and3_1
XANTENNA__09532__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08429__B net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08584_ net781 net766 _04715_ net681 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14252__A2 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12666__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1081_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout437_A _08022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17316__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1179_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\] net658 net609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\]
+ _05451_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout604_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ net1075 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] net873
+ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__and3_1
XANTENNA__17466__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[18\] net910
+ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__and3_1
XANTENNA__15278__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold650 team_01_WB.instance_to_wrap.cpu.f0.num\[14\] vssd1 vssd1 vccd1 vccd1 net2266
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09707__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\] vssd1 vssd1 vccd1 vccd1 net2288
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _03392_ vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16490__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold694 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13279__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] net657 net632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11829__A1 _07551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ net1885 net605 net587 _03661_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a22o_1
Xhold1350 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1361 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2977 sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ net2565 net291 net476 vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1372 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14650_ net1404 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
X_11862_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[7\] net677 net778 vssd1 vssd1
+ vccd1 vccd1 _07979_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14243__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ net768 _07265_ net1066 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__o21a_1
X_10813_ _07073_ _07075_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__nand2_1
X_14581_ net1205 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XANTENNA__12576__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ _07858_ _07921_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__or2_1
X_16320_ clknet_leaf_75_wb_clk_i net1965 _00188_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13532_ _07881_ _03881_ net185 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10744_ _05852_ _05788_ net504 vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17809__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16251_ clknet_leaf_69_wb_clk_i _01888_ _00119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13463_ _03814_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__and2_1
X_10675_ _06664_ _06643_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_129_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15202_ net1266 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12414_ net1978 net250 net421 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
X_16182_ clknet_leaf_90_wb_clk_i _01850_ _00050_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11216__A_N _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13394_ net2619 net327 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1
+ vccd1 vccd1 _01889_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15133_ net1283 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ net3085 net219 net490 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08630__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13200__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09186__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15064_ net1254 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XANTENNA__08090__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12276_ net2562 net229 net431 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03577_ _04142_ _00005_ vssd1
+ vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_read_i sky130_fd_sc_hd__a31o_1
X_11227_ net321 _07486_ _07490_ _07106_ _07489_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__a221o_1
XANTENNA__10125__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09914__A _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ _06319_ _06887_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__or2_1
XANTENNA__16983__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\] _04774_ _06352_
+ _06359_ _06368_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__a2111o_1
X_15966_ net1336 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__inv_2
X_11089_ _06110_ net342 net335 _06108_ net333 vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__a221o_1
X_14917_ net1225 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
X_17705_ clknet_leaf_110_wb_clk_i _03265_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12493__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ net1350 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__inv_2
XANTENNA__17339__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17636_ clknet_leaf_138_wb_clk_i _03196_ _01499_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14848_ net1359 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12486__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17567_ clknet_leaf_1_wb_clk_i _03127_ _01430_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08449__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12245__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ net1407 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ clknet_leaf_73_wb_clk_i _02146_ _00381_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10256__B1 _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17498_ clknet_leaf_36_wb_clk_i _03058_ _01361_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16363__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18231__1590 vssd1 vssd1 vccd1 vccd1 _18231__1590/HI net1590 sky130_fd_sc_hd__conb_1
XFILLER_0_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11403__B _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16449_ clknet_leaf_98_wb_clk_i _02077_ _00312_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09413__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18119_ net1493 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08621__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13110__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09096__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__C _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15826__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout404 _03563_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_4
XANTENNA__10035__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout415 net418 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_8
Xfanout426 _08027_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout437 _08022_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_8
X_09823_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] net879 vssd1
+ vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__and3_1
XANTENNA__09824__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout448 _08019_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_4
Xfanout459 _08015_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_6
XFILLER_0_96_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] net610 _06002_
+ _06003_ _06007_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_119_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] net920 vssd1
+ vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__and3_1
X_09685_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\] net636 _05925_
+ _05930_ _05934_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08688__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09262__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1296_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08636_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] _04741_ net613
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] _04889_ vssd1 vssd1 vccd1
+ vccd1 _04900_ sky130_fd_sc_hd__a221o_1
XANTENNA__10201__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16706__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12396__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] net664 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout721_A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout819_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08498_ net1068 net896 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__and2_2
XFILLER_0_119_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10262__A3 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\] net730 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09119_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] net898
+ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__and3_1
XANTENNA__08612__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ _06648_ _06650_ _06652_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12130_ net2162 net309 net454 vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__mux2_1
XANTENNA__09437__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ net2643 net260 net461 vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\] vssd1 vssd1 vccd1 vccd1
+ net2096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold491 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[3\] vssd1 vssd1 vccd1 vccd1
+ net2107 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__A3 _07734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ _07027_ _07031_ net513 vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15820_ net1252 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__inv_2
Xfanout971 net973 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 _04485_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15751_ net1184 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
X_12963_ net1033 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\] vssd1 vssd1 vccd1
+ vccd1 _03649_ sky130_fd_sc_hd__or2_1
XANTENNA__08679__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1180 team_01_WB.instance_to_wrap.cpu.f0.num\[7\] vssd1 vssd1 vccd1 vccd1 net2796
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08143__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14702_ net1377 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
X_11914_ net2386 net254 net476 vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15682_ net1267 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ net1025 _07653_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ clknet_leaf_21_wb_clk_i _02981_ _01284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14633_ net1386 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XANTENNA__17631__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\] net679 net780 vssd1 vssd1
+ vccd1 vccd1 _07965_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17352_ clknet_leaf_45_wb_clk_i _02912_ _01215_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14564_ net1324 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ _07860_ _07907_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16303_ clknet_leaf_113_wb_clk_i _01937_ _00171_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] _04727_ vssd1 vssd1
+ vccd1 vccd1 _03868_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11223__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17283_ clknet_leaf_119_wb_clk_i _02843_ _01146_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ _06845_ _06952_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__or2_4
X_14495_ net1339 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17781__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16234_ clknet_leaf_38_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[15\]
+ _00102_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18096__1470 vssd1 vssd1 vccd1 vccd1 _18096__1470/HI net1470 sky130_fd_sc_hd__conb_1
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13446_ _03797_ _03798_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__or2_1
X_10658_ _06919_ _06921_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__and2_1
XANTENNA__08813__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16165_ clknet_leaf_57_wb_clk_i _01833_ _00033_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08603__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13377_ net2324 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1
+ vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
X_10589_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _06847_ _04725_ vssd1 vssd1
+ vccd1 vccd1 _06853_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ net1263 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
X_12328_ net2306 net308 net430 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XANTENNA__12950__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16096_ net1376 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15047_ net1181 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
X_12259_ net2023 net298 net438 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17161__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16998_ clknet_leaf_140_wb_clk_i _02558_ _00861_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15949_ net1393 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15381__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] net850
+ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__and3_1
XANTENNA__14207__A2 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10021__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ net980 net950 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17619_ clknet_leaf_21_wb_clk_i _03179_ _01482_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09810__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16879__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\] net3241 net1042 vssd1 vssd1
+ vccd1 vccd1 _03395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08283_ net3181 net3160 net1049 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_138_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09819__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout302_A _07970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10691__C _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09257__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16259__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17504__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1211_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 _07906_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout212 net214 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1309_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout223 _07915_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xfanout234 net237 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
XANTENNA_fanout671_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 _07980_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xfanout256 net258 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_2
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 net269 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
X_09806_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] net710 net758 vssd1
+ vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__o21ai_1
Xfanout278 net281 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
XANTENNA_hold1417_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__A2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 _07901_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] net872
+ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__and3_1
XANTENNA__17654__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09668_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\] net894 vssd1
+ vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__and3_1
XANTENNA__09873__A2 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] net759 _04881_ _04882_
+ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a22o_2
X_09599_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] net878 vssd1
+ vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__and3_1
XANTENNA__13015__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11630_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[11\] _07806_ vssd1 vssd1 vccd1
+ vccd1 _07830_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A2 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _04478_ _07731_ _07770_ _07789_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a31o_1
XANTENNA__12854__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13300_ net1758 net808 net803 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\] vssd1
+ vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13709__A1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10512_ _06752_ _06774_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17034__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14280_ _04158_ _04288_ _04413_ _04433_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__nor4_1
X_11492_ _07731_ _07740_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09389__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13231_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] net3244 net831 vssd1 vssd1
+ vccd1 vccd1 _02027_ sky130_fd_sc_hd__mux2_1
X_10443_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\] net646 net616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__a22o_1
XANTENNA__11196__B2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input65_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ net2202 net1956 net818 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09167__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _06624_ _06635_ _06636_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10943__A1 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12113_ net2336 net285 net451 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__mux2_1
X_13093_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\] net1028 vssd1 vssd1 vccd1
+ vccd1 _03716_ sky130_fd_sc_hd__or2_1
X_17970_ clknet_leaf_89_wb_clk_i _03519_ _01790_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.read_i
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09464__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ net2226 net226 net459 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
X_16921_ clknet_leaf_17_wb_clk_i _02481_ _00784_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16852_ clknet_leaf_7_wb_clk_i _02412_ _00715_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout790 _04228_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_2
X_15803_ net1297 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16783_ clknet_leaf_54_wb_clk_i _02343_ _00646_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13995_ _03554_ _03553_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15734_ net1304 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12946_ net1027 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[11\] vssd1 vssd1 vccd1
+ vccd1 _03637_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11120__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09864__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11120__B2 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15665_ net1189 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XANTENNA__09630__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] net1056 net366 _03586_
+ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14616_ net1406 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17404_ clknet_leaf_14_wb_clk_i _02964_ _01267_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11828_ net780 _07950_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15596_ net1265 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09616__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17335_ clknet_leaf_9_wb_clk_i _02895_ _01198_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14547_ net1324 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11759_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _07861_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12764__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08824__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17266_ clknet_leaf_39_wb_clk_i _02826_ _01129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09639__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14478_ net1392 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08543__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16217_ clknet_leaf_116_wb_clk_i _01884_ _00085_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13429_ _03780_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17197_ clknet_leaf_16_wb_clk_i _02757_ _01060_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16148_ net1338 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_max_cap901_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] net733 net716 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ net1368 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_100_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14280__A _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10016__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17677__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10698__A0 _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XFILLER_0_78_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _05778_ _05779_ _05784_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] net710 net758 vssd1
+ vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__o21a_1
XANTENNA__09540__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout252_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08404_ net1147 net1152 net1154 net1149 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09384_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\] net735 net711 _05646_
+ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_47_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08335_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12674__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14455__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1259_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ net2259 net2058 net1047 vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08197_ _04554_ _04583_ _04587_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout886_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1007 net1008 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
X_10090_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\] net874 vssd1
+ vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1018 net1023 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_2
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_105_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12849__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12800_ net3210 net204 net373 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13780_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] _04084_ _04085_ vssd1 vssd1 vccd1
+ vccd1 _04086_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_74_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ net530 _07182_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13948__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10877__B _07140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ net3057 net190 net379 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15450_ net1260 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
X_12662_ net2972 net213 net394 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ net1351 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
X_11613_ net496 _07821_ net2096 net839 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__o2bb2a_1
X_15381_ net1178 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
XANTENNA__12584__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ net2155 net307 net402 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
XANTENNA__16424__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ clknet_leaf_142_wb_clk_i _02680_ _00983_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1
+ vccd1 _02266_ sky130_fd_sc_hd__clkbuf_1
X_11544_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] _07777_ vssd1 vssd1 vccd1 vccd1
+ _07779_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09459__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__A team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ clknet_leaf_32_wb_clk_i _02611_ _00914_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\] _04267_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\]
+ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a221o_1
X_11475_ _04462_ _04505_ _07727_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__or3b_1
XFILLER_0_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16002_ net1394 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__inv_2
XANTENNA__11169__B2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13214_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\]
+ net821 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10426_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\] net731 net724 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__a22o_1
XANTENNA__16574__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194_ net147 net585 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11928__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ net2347 net1633 net828 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__mux2_1
X_10357_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\] net914
+ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10392__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ _06105_ _07806_ net1026 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__o21a_1
XANTENNA__13428__B _06348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17953_ clknet_leaf_107_wb_clk_i _03503_ _01773_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10288_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\] net853 vssd1
+ vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16904_ clknet_leaf_63_wb_clk_i _02464_ _00767_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12027_ net3139 net300 net465 vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
X_17884_ clknet_leaf_75_wb_clk_i _03434_ _01704_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11341__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09922__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16835_ clknet_leaf_131_wb_clk_i _02395_ _00698_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12759__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13094__A1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13978_ _04167_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__inv_2
X_16766_ clknet_leaf_13_wb_clk_i _02326_ _00629_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08538__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15717_ net1225 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
X_12929_ team_01_WB.instance_to_wrap.a1.ADR_I\[16\] net604 net586 _03624_ vssd1 vssd1
+ vccd1 vccd1 _02224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12841__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16697_ clknet_leaf_123_wb_clk_i _02257_ _00560_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09360__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ net1276 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15579_ net1318 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
XANTENNA__12494__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ _04531_ _04532_ _04546_ _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__and4b_1
XFILLER_0_71_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17318_ clknet_leaf_139_wb_clk_i _02878_ _01181_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09369__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08704__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17249_ clknet_leaf_136_wb_clk_i _02809_ _01112_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10308__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08576__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10383__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08953_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\] net937
+ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09535__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15834__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08884_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] net918 vssd1
+ vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1007_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__B2 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12669__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18075__1449 vssd1 vssd1 vccd1 vccd1 _18075__1449/HI net1449 sky130_fd_sc_hd__conb_1
XANTENNA__13085__A1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11096__A0 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09505_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\] net922 vssd1
+ vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09270__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11635__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1376_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09436_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] net944
+ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13801__B team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09367_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[13\] net961
+ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__and3_1
XANTENNA__14185__A _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ net2679 net2640 net1041 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
X_09298_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\] net930
+ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17842__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08249_ net2480 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ _05622_ _06907_ _07200_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__and3b_1
XANTENNA__09213__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12899__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08911__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\] net740 net723 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__a22o_1
XANTENNA__08567__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ net547 _07452_ _07454_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10142_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\] net703 _06387_ _06388_
+ _06395_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__a2111o_1
X_10073_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\] _04648_ net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[3\]
+ _06332_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__a221o_1
X_14950_ net1281 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XANTENNA__09742__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] net795 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[14\] sky130_fd_sc_hd__and2_1
X_14881_ net1314 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12579__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13832_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[4\] team_01_WB.instance_to_wrap.cpu.c0.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__and4bb_1
X_16620_ clknet_leaf_86_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[6\]
+ _00483_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13076__A1 _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16551_ clknet_leaf_47_wb_clk_i _02179_ _00414_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ _04470_ _04072_ _04015_ _04558_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_74_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12823__A1 _07994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10975_ _07137_ _07144_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__a21oi_1
X_15502_ net1217 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
X_12714_ net2921 net274 net384 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16482_ clknet_leaf_108_wb_clk_i _02110_ _00345_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_13694_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _04015_ vssd1 vssd1 vccd1 vccd1
+ _04016_ sky130_fd_sc_hd__nand2_1
XANTENNA__11215__C _07456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15433_ net1214 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
X_18221_ net601 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_1
X_12645_ net2180 net250 net393 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XANTENNA__10827__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10047__D1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11512__A team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18152_ net1526 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XFILLER_0_93_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15364_ net1226 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XANTENNA__09189__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__A team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12576_ net2094 net283 net401 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17103_ clknet_leaf_19_wb_clk_i _02663_ _00966_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14315_ net1366 _04453_ _04454_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nor3_1
X_11527_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] _07745_ _07762_ _07764_ vssd1
+ vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__o211a_1
X_18083_ net1457 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15295_ net1295 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10128__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ clknet_leaf_41_wb_clk_i _02594_ _00897_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold309 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] _04238_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\]
+ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11458_ _04471_ _07710_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\] net929
+ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14177_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\] _04242_ _04280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\]
+ _04335_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ net344 _07641_ _07647_ _07652_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13128_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\] net2775 net827 vssd1 vssd1
+ vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13059_ net1971 net834 net355 _03692_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17936_ clknet_leaf_101_wb_clk_i _03486_ _01756_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1009 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1360 net1414 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__clkbuf_2
Xfanout1371 net1379 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__buf_4
Xfanout1382 net1389 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__buf_4
X_17867_ clknet_leaf_80_wb_clk_i net2687 _01687_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12489__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1393 net1398 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08730__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16818_ clknet_leaf_31_wb_clk_i _02378_ _00681_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17798_ clknet_leaf_69_wb_clk_i _03355_ _01619_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16749_ clknet_leaf_21_wb_clk_i _02309_ _00612_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09090__C _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10825__A0 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13902__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _05482_ _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__or2_2
XFILLER_0_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _05415_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__inv_2
XANTENNA__09443__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _04496_ team_01_WB.instance_to_wrap.cpu.f0.num\[8\]
+ _04477_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__o22a_1
XANTENNA__08797__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15829__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _05309_ _05345_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__nand2_2
XANTENNA__10038__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _07943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08034_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 _04465_
+ sky130_fd_sc_hd__inv_2
Xinput70 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09827__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold810 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold821 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold832 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 team_01_WB.instance_to_wrap.cpu.c0.count\[16\] vssd1 vssd1 vccd1 vccd1 net2459
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11002__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold854 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[26\] vssd1 vssd1 vccd1 vccd1
+ net2470 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold865 _03498_ vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold876 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13068__B net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17245__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\] net918 vssd1
+ vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__and3_1
XANTENNA__09265__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout584_A _04157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ net583 _05167_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__or2_1
XANTENNA__10108__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10204__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1510 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09562__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1532 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3148 sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[20\] net608 _05103_
+ _05104_ _05106_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout751_A _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1543 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] vssd1 vssd1 vccd1 vccd1
+ net3181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17395__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1576 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3192 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08721__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1587 team_01_WB.instance_to_wrap.cpu.f0.num\[3\] vssd1 vssd1 vccd1 vccd1 net3203
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08798_ _05057_ _05058_ _05059_ _05061_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nor4_1
Xhold1598 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10760_ _04854_ _06841_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08906__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09419_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\] net609 _05655_
+ _05659_ _05664_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10691_ net542 net538 _06953_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__and3_2
X_12430_ net2068 net290 net420 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12361_ net3169 net309 net493 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11241__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14100_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[112\] _04260_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\]
+ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__a22o_1
XANTENNA__11792__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ _06963_ _07007_ net526 vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09737__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15080_ net1208 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
X_12292_ net3201 net300 net434 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14031_ _04509_ _04146_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nand2_1
XANTENNA__13259__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11243_ net321 _07140_ _07503_ _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11174_ _07405_ _07407_ net529 vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10125_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\] net952 vssd1
+ vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__and3_1
XANTENNA__15474__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16612__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15982_ net1386 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__inv_2
X_17721_ clknet_leaf_110_wb_clk_i _03281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09472__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] net925 vssd1
+ vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14933_ net1177 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08712__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12102__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17652_ clknet_leaf_4_wb_clk_i _03212_ _01515_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08088__A team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10411__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ net1346 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XANTENNA__14246__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16603_ clknet_leaf_118_wb_clk_i _02231_ _00466_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13815_ net2146 net785 _04559_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1
+ vccd1 vccd1 _01827_ sky130_fd_sc_hd__a22o_1
X_14795_ net1334 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17583_ clknet_leaf_18_wb_clk_i _03143_ _01446_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11941__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16534_ clknet_leaf_60_wb_clk_i _02162_ _00397_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13746_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] net783 _04057_ _04059_
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10958_ net345 _07220_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08816__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13441__B net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13677_ _03782_ _03786_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__xor2_1
XANTENNA__17118__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16465_ clknet_leaf_99_wb_clk_i _02093_ _00328_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10889_ net344 _07125_ _07130_ _07151_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ net1578 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
X_12628_ net2380 net290 net397 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
X_15416_ net1257 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
X_16396_ clknet_leaf_101_wb_clk_i _02024_ _00259_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18135_ net1509 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
X_15347_ net1178 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XANTENNA__08779__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ net2067 net313 net405 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__mux2_1
XANTENNA__12772__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12980__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18066_ net1440 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15278_ net1214 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
Xhold106 _03514_ vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18074__1448 vssd1 vssd1 vccd1 vccd1 _18074__1448/HI net1448 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold117 _02063_ vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\] vssd1 vssd1 vccd1 vccd1
+ net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 team_01_WB.instance_to_wrap.cpu.f0.write_data\[7\] vssd1 vssd1 vccd1 vccd1
+ net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13524__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17017_ clknet_leaf_18_wb_clk_i _02577_ _00880_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14229_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\] _04255_ _04272_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\]
+ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout619 _04771_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15384__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09770_ _05761_ _06033_ _05756_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__o21a_1
XANTENNA__10024__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] net753 net711 _04965_
+ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a2111o_1
X_17919_ clknet_leaf_108_wb_clk_i net2131 _01739_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1190 net1194 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08652_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] net913 vssd1
+ vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__and3_1
XANTENNA__12012__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ _04832_ _04833_ _04846_ net666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__o32a_4
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11851__S net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout332_A _06989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1074_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09204_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\] net640 _05452_ _05455_
+ _05458_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09135_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\] net908
+ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12682__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14463__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1339_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12971__B1 _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\] net903
+ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08461__A team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14182__B _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout799_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16635__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold651 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold673 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\] net661 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__a22o_1
XANTENNA__09292__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16785__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] net873 vssd1
+ vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] net665 _06152_ _06157_
+ _06158_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__a2111o_1
Xhold1340 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13018__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ net2097 net295 net478 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_1
Xhold1351 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10231__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1362 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13245__C net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1373 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14228__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1384 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1395 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11861_ net677 _07368_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__nand2_1
XANTENNA__12857__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11761__S net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ net768 _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__nand2_1
XANTENNA__13542__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10812_ net542 _07074_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14580_ net1344 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09655__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _07857_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\]
+ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _03757_ _03864_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _07005_ _07006_ net516 vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16250_ clknet_leaf_70_wb_clk_i _01887_ _00118_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13462_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _05584_ vssd1 vssd1
+ vccd1 vccd1 _03815_ sky130_fd_sc_hd__xor2_1
X_10674_ _06752_ _06775_ _06937_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15201_ net1291 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12413_ net2318 net254 net420 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XANTENNA__15469__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16181_ clknet_leaf_90_wb_clk_i _01849_ _00049_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12592__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ net2375 net329 net353 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1
+ vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14373__A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15132_ net1232 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09467__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ net2458 net284 net492 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08371__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10973__C1 _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ net1250 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09186__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12275_ net3062 net200 net431 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10406__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11517__A1 _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03581_ _04142_ vssd1 vssd1
+ vccd1 vccd1 _00006_ sky130_fd_sc_hd__and3_1
X_11226_ _07249_ _07438_ net535 vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11936__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ net547 _07415_ _07420_ _07106_ _07418_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10108_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[3\] net619 _06361_ _06363_
+ _06369_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15965_ net1336 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__inv_2
XANTENNA__09633__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11088_ _06967_ _07211_ net531 vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17704_ clknet_leaf_110_wb_clk_i _03264_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10039_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] net639 _06281_ _06297_
+ _06301_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a2111o_1
X_14916_ net1269 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XANTENNA__14219__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15896_ net1354 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__inv_2
XANTENNA__09930__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17635_ clknet_leaf_119_wb_clk_i _03195_ _01498_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14847_ net1384 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XANTENNA__12767__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_125_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17566_ clknet_leaf_13_wb_clk_i _03126_ _01429_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14778_ net1334 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XANTENNA__09646__B1 _04685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08546__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16508__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09110__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16517_ clknet_leaf_72_wb_clk_i _02145_ _00380_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13729_ _04026_ _04046_ net485 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17497_ clknet_leaf_17_wb_clk_i _03057_ _01360_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16448_ clknet_leaf_106_wb_clk_i _02076_ _00311_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16379_ clknet_leaf_112_wb_clk_i net1750 _00247_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10559__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11700__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12953__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18118_ net1492 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
XANTENNA__17903__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18049_ net1611 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_83_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12007__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09177__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14170__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout405 _03563_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_8
Xfanout416 net418 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_4
X_09822_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] net852 vssd1
+ vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__and3_1
Xfanout427 _08024_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08924__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13627__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10750__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _08022_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout449 _08019_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_8
X_09753_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] net660 _05996_ _06005_
+ _06010_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09543__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_A _07920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] net950 vssd1
+ vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__and3_1
X_09684_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\] net617 _05933_ _05940_
+ _05942_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13681__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08635_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\] net657 _04898_
+ net672 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a211o_1
XANTENNA__12677__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14458__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A _06314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1191_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1289_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\] net637 net612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18189__1563 vssd1 vssd1 vccd1 vccd1 _18189__1563/HI net1563 sky130_fd_sc_hd__conb_1
XANTENNA__09101__A2 _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08497_ net1081 net851 vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__and2_2
XFILLER_0_18_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17583__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12944__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ net1075 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] net905
+ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10390_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\] net628 net621 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\]
+ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09049_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] net845
+ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14921__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ net2217 net299 net462 vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14161__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold470 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net330 _06995_ _07272_ net540 _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout950 net952 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_4
Xfanout961 net964 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_8
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout983 net992 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net1009 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ net1293 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
X_12962_ net1033 _07396_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__nand2_1
Xhold1170 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 net2786
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net2439 net220 net476 vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\] vssd1 vssd1 vccd1 vccd1
+ net2797 sky130_fd_sc_hd__dlygate4sd3_1
X_14701_ net1375 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1192 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 net2808
+ sky130_fd_sc_hd__dlygate4sd3_1
X_15681_ net1292 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XANTENNA__12587__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ net1953 net607 net589 _03598_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
X_18073__1447 vssd1 vssd1 vccd1 vccd1 _18073__1447/HI net1447 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17420_ clknet_leaf_44_wb_clk_i _02980_ _01283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ net1406 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
X_11844_ _07852_ _07963_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ net1322 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_17351_ clknet_leaf_121_wb_clk_i _02911_ _01214_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13975__A2 _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07859_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\]
+ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__a21oi_1
X_16302_ clknet_leaf_112_wb_clk_i _01936_ _00170_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16800__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13514_ _03753_ _03866_ _03752_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21bo_1
X_10726_ _06845_ _06952_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__nor2_1
XANTENNA__17926__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ net1343 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
X_17282_ clknet_leaf_142_wb_clk_i _02842_ _01145_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16233_ clknet_leaf_37_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[14\]
+ _00101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13445_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _05924_ _03794_ _03795_
+ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__nor4_1
X_10657_ _05419_ _05486_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11520__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09197__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ net3155 net328 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1
+ vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
X_16164_ clknet_leaf_90_wb_clk_i _01832_ _00032_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10588_ _04726_ _06851_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__nor2_1
XANTENNA__09800__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16950__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12327_ net2292 net312 net430 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
X_15115_ net1221 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
X_16095_ net1366 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15046_ net1274 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14152__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ net2368 net242 net436 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
XANTENNA__13447__A team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11209_ net537 _07069_ _07472_ _07471_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__a31o_1
XANTENNA__13360__B1 _03747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17306__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ net3171 net265 net444 vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09363__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16997_ clknet_leaf_131_wb_clk_i _02557_ _00860_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15948_ net1391 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10302__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12497__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15879_ net1356 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08420_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\] net914 vssd1
+ vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17618_ clknet_leaf_22_wb_clk_i _03178_ _01481_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] net1826 net1047 vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08707__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17549_ clknet_leaf_19_wb_clk_i _03109_ _01412_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16480__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ net2019 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\] net1052 vssd1 vssd1
+ vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09538__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15837__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1037_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10952__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14143__A2 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12154__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13351__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _07888_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
XFILLER_0_10_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout224 _07915_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
Xfanout235 net237 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_1
X_09805_ _06058_ _06063_ _06066_ _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__nor4_1
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
Xfanout279 net281 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09273__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\] net903
+ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09570__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\] net862
+ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and3_1
XANTENNA__11665__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout831_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout929_A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17949__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\] net846 vssd1
+ vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__and3_1
XANTENNA__11417__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] net729 _04801_
+ _04806_ _04807_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ net320 _07788_ net1065 vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08914__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16973__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10511_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11491_ _07721_ _07739_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ net823 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10442_ _06699_ _06701_ _06703_ _06705_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11196__A2 _06983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__A1 _07989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13966__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ net3004 net2862 net828 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13590__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10373_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] net743 net706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10943__A2 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ net2267 net225 net452 vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__mux2_1
XANTENNA__09745__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14134__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input58_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _05820_ _07807_ _03704_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13342__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16920_ clknet_leaf_23_wb_clk_i _02480_ _00783_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12043_ net1927 net200 net459 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XANTENNA__16353__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16851_ clknet_leaf_49_wb_clk_i _02411_ _00714_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout780 _04623_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout791 _04224_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__buf_2
X_15802_ net1257 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16782_ clknet_leaf_53_wb_clk_i _02342_ _00645_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13994_ _04163_ _03553_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09313__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15733_ net1179 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ net1027 _07568_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08521__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13206__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12110__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15664_ net1247 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
X_12876_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] _07082_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17403_ clknet_leaf_32_wb_clk_i _02963_ _01266_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14615_ net1372 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
X_11827_ _07854_ _07949_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__or2_1
X_15595_ net1210 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XANTENNA__11959__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13730__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17334_ clknet_leaf_29_wb_clk_i _02894_ _01197_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14546_ net1317 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
X_11758_ net2485 net237 net479 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18019__1596 vssd1 vssd1 vccd1 vccd1 net1596 _18019__1596/LO sky130_fd_sc_hd__conb_1
XFILLER_0_43_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10709_ _06807_ _06752_ net498 vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__mux2_1
X_17265_ clknet_leaf_21_wb_clk_i _02825_ _01128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ net2792 _07837_ net35 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a21o_1
X_14477_ net1392 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16216_ clknet_leaf_117_wb_clk_i _01883_ _00084_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_13428_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _06348_ vssd1 vssd1 vccd1
+ vccd1 _03781_ sky130_fd_sc_hd__or2_1
X_17196_ clknet_leaf_46_wb_clk_i _02756_ _01059_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13581__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16147_ net1325 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12780__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ net28 net800 net595 net1846 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10395__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14125__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ net1372 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13333__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15029_ net1173 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10147__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18188__1562 vssd1 vssd1 vccd1 vccd1 _18188__1562/HI net1562 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09552__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A1 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09093__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13905__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10032__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[9\] net726 net712 _05768_
+ _05773_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09390__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09821__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11425__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _05706_ _05708_ _05712_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__or4_4
XANTENNA__12020__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08403_ net1117 net928 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and2_4
XANTENNA__16996__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09383_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] net748 _05624_
+ _05629_ _05633_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout245_A _07980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08334_ net2552 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\] net1041 vssd1 vssd1
+ vccd1 vccd1 _03413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\] net1791 net1050 vssd1 vssd1
+ vccd1 vccd1 _03482_ sky130_fd_sc_hd__mux2_1
XANTENNA__10622__B2 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout412_A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1154_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ net1813 net553 _04568_ _04595_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09268__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12690__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1321_A net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10386__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18072__1446 vssd1 vssd1 vccd1 vccd1 _18072__1446/HI net1446 sky130_fd_sc_hd__conb_1
XFILLER_0_105_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09565__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout781_A _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13324__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_A _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1019 net1022 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08909__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09719_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] net741 _05966_ _05971_
+ _05975_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09731__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ _05417_ net337 _07254_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_134_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12730_ net1938 net196 net380 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XANTENNA__13253__C _03734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17001__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ net2906 net291 net392 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[20\] net573 vssd1 vssd1 vccd1
+ vccd1 _07821_ sky130_fd_sc_hd__nand2_1
X_14400_ net1352 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12592_ net3211 net311 net402 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__mux2_1
X_15380_ net1243 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08644__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ net483 _07777_ net319 vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ net2103 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08363__B net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17050_ clknet_leaf_32_wb_clk_i _02610_ _00913_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] _04242_ _04275_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\]
+ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a22o_1
X_11474_ _07721_ _07724_ _07726_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__and3_1
XANTENNA__16719__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16001_ net1363 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10425_ _06685_ _06686_ _06687_ _06688_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__or4_1
XANTENNA__15477__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14193_ _04330_ _04339_ _04345_ _04351_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13144_ net2797 net1640 net827 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
X_10356_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\] net958
+ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08810__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13075_ net3046 net835 net354 _03703_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
X_17952_ clknet_leaf_100_wb_clk_i _03502_ _01772_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[0\] net844 vssd1
+ vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__and3_1
XANTENNA__10414__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12105__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12332__C _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13866__B2 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16903_ clknet_leaf_133_wb_clk_i _02463_ _00766_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12026_ net2716 net244 net465 vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
X_17883_ clknet_leaf_80_wb_clk_i _03433_ _01703_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08742__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11944__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16834_ clknet_leaf_144_wb_clk_i _02394_ _00697_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08819__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16765_ clknet_leaf_129_wb_clk_i _02325_ _00628_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09641__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ net1170 _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__nand2_2
XFILLER_0_92_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15716_ net1270 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
X_12928_ net364 _03622_ _03623_ net1053 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a32o_1
X_16696_ clknet_leaf_25_wb_clk_i _02256_ _00559_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10793__A2_N net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15647_ net1295 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XANTENNA__12775__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16249__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ net2409 net290 net369 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11899__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15578_ net1305 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17317_ clknet_leaf_133_wb_clk_i _02877_ _01180_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14529_ net1323 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16399__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 _04481_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10080__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17248_ clknet_leaf_142_wb_clk_i _02808_ _01111_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09088__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09758__C1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17179_ clknet_leaf_39_wb_clk_i _02739_ _01042_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10368__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10027__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09816__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13306__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12015__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] net950 vssd1
+ vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__and3_1
XANTENNA__17794__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\] net958 vssd1
+ vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and3_1
XANTENNA__08733__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17024__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout362_A _03665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09504_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\] _04641_ net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a22o_1
XANTENNA__11096__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09435_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\] net917
+ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12685__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14466__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17174__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1271_A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout627_A _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1369_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09366_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] net940
+ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14185__B _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08317_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] net2358 net1044 vssd1 vssd1
+ vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] net941
+ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__and3_1
XANTENNA_hold1477_A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10071__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout996_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08179_ _04553_ _04572_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12899__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] net705 net695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ _06473_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09295__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _07118_ _07237_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08972__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\] net690 _06391_ _06393_
+ _06396_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__a2111o_1
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_101_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09516__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _06329_ _06333_ _06334_ _06335_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11859__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__B1 _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18018__1595 vssd1 vssd1 vccd1 vccd1 net1595 _18018__1595/LO sky130_fd_sc_hd__conb_1
X_13900_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] net797 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[13\] sky130_fd_sc_hd__and2_1
X_14880_ net1311 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
XANTENNA__10531__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ _04122_ _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nor2_1
XANTENNA__09461__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13076__A2 _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17517__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16550_ clknet_leaf_41_wb_clk_i _02178_ _00413_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13762_ _07713_ _07773_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nand2_1
X_10974_ _06970_ _07143_ _07237_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15501_ net1213 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ net2363 net218 net384 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XANTENNA__12595__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16481_ clknet_leaf_99_wb_clk_i _02109_ _00344_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_112_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13693_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] net1063 team_01_WB.instance_to_wrap.cpu.f0.i\[16\]
+ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__and4_1
X_18220_ net602 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_1
X_15432_ net1185 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
X_12644_ net3247 net257 net392 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18187__1561 vssd1 vssd1 vccd1 vccd1 _18187__1561/HI net1561 sky130_fd_sc_hd__conb_1
XFILLER_0_66_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18151_ net1525 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12575_ net2892 net224 net401 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15363_ net1219 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10409__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ clknet_leaf_55_wb_clk_i _02662_ _00965_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14314_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ _04450_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and3_1
X_11526_ _04471_ _07710_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__nand2_1
X_18082_ net1456 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XFILLER_0_81_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15294_ net1316 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17033_ clknet_leaf_40_wb_clk_i _02593_ _00896_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11939__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07708_ vssd1 vssd1 vccd1 vccd1
+ _07710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14245_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\] _04242_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10408_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\] net929 vssd1
+ vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09755__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14176_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\] _04233_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[43\]
+ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a22o_1
XANTENNA__11011__B2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ _07080_ _07648_ _07651_ _07643_ _07646_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09636__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08540__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__A2 _07734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13127_ net3048 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\] net831 vssd1 vssd1
+ vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
X_10339_ _06180_ _06319_ _06597_ _06600_ _06177_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__o41a_2
XANTENNA__10770__A0 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17047__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[20\] _03691_ net1028 vssd1
+ vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__mux2_1
XANTENNA__09507__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17935_ clknet_leaf_109_wb_clk_i net2788 _01755_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12511__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08715__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ net2270 net288 net463 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__mux2_1
Xfanout1350 net1351 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__buf_4
XANTENNA__13455__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1361 net1362 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__buf_4
X_17866_ clknet_leaf_78_wb_clk_i _03416_ _01686_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1372 net1379 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__clkbuf_4
Xfanout1383 net1389 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1394 net1395 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__buf_4
XFILLER_0_89_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16817_ clknet_leaf_21_wb_clk_i _02377_ _00680_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_17797_ clknet_leaf_70_wb_clk_i _03354_ _01618_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15670__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16748_ clknet_leaf_45_wb_clk_i _02308_ _00611_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10310__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10825__A1 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18071__1445 vssd1 vssd1 vccd1 vccd1 _18071__1445/HI net1445 sky130_fd_sc_hd__conb_1
XANTENNA__13902__B net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16679_ clknet_leaf_105_wb_clk_i net795 _00542_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.ihit
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _05448_ _05481_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11703__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09151_ _05379_ _05414_ net583 vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_2
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _04491_ _04493_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09082_ _05309_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__nor2_1
XANTENNA__11250__B2 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 _04464_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_13_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold800 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xinput60 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xhold811 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] vssd1 vssd1 vccd1 vccd1
+ net2427 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout208_A _07879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold822 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold833 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13938__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold844 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\] vssd1 vssd1 vccd1 vccd1
+ net2482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold877 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\] vssd1 vssd1 vccd1 vccd1
+ net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\] net915 vssd1
+ vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__and3_1
Xhold899 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1117_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08935_ _05195_ _05197_ _05198_ _05168_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__o31a_4
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1500 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[0\] vssd1 vssd1 vccd1 vccd1
+ net3116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3149 sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\] _04749_ _05105_
+ _05108_ _05121_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a2111o_1
Xhold1544 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\] vssd1 vssd1 vccd1 vccd1
+ net3160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08459__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1555 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1566 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 team_01_WB.instance_to_wrap.cpu.f0.num\[25\] vssd1 vssd1 vccd1 vccd1 net3193
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08797_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\] net662 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\]
+ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout744_A _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1588 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1599 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16564__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\] net617 _05681_ net671
+ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a211oi_1
X_10690_ net542 _06953_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13766__B1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09349_ _05609_ _05610_ _05611_ _05612_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10044__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12360_ net2920 net313 net493 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08922__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13518__A0 _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11311_ _07004_ _07555_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__nand2_1
X_12291_ net2294 net242 net433 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__mux2_1
X_14030_ _04146_ net565 _04204_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__and3_1
XANTENNA__14191__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ _06030_ net341 _07505_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13259__B net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12741__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ net523 _07404_ net535 vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10752__A0 _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input40_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] net952 vssd1
+ vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15981_ net1386 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17720_ clknet_leaf_110_wb_clk_i _03280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10055_ _06316_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__nand2_2
X_14932_ net1238 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XANTENNA__10504__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17651_ clknet_leaf_50_wb_clk_i _03211_ _01514_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14863_ net1341 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ clknet_leaf_78_wb_clk_i _02230_ _00465_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13814_ net2009 net785 _04559_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1
+ vccd1 vccd1 _01828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17582_ clknet_leaf_55_wb_clk_i _03142_ _01445_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ net1328 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10130__C _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16533_ clknet_leaf_67_wb_clk_i _02161_ _00396_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ net485 _04058_ net785 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a21o_1
X_10957_ _05621_ _07205_ _06036_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13214__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10283__A2 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ clknet_leaf_106_wb_clk_i _02092_ _00327_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13676_ net968 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _04000_ _04001_
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10888_ net344 _07125_ _07130_ _07151_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18203_ net1577 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XFILLER_0_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15415_ net1250 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
X_12627_ net2706 net296 net398 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16395_ clknet_leaf_76_wb_clk_i _02023_ _00258_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08228__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18134_ net1508 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
XFILLER_0_109_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15346_ net1174 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12558_ net2243 net259 net406 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11783__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12980__B2 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18065_ net1439 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
X_11509_ team_01_WB.instance_to_wrap.cpu.f0.i\[22\] _07745_ _07750_ _07752_ vssd1
+ vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ net1213 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
Xhold107 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 net1723
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ net2826 net316 net412 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 team_01_WB.instance_to_wrap.a1.ADR_I\[14\] vssd1 vssd1 vccd1 vccd1 net1734
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17016_ clknet_leaf_27_wb_clk_i _02576_ _00879_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold129 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\] vssd1 vssd1 vccd1 vccd1
+ net1745 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\] _04266_ _04280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\]
+ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09366__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14159_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\] _04261_ _04280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[98\]
+ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__a221o_1
Xfanout609 _04777_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_6
XANTENNA__10305__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08720_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] net742 _04963_
+ _04967_ _04971_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17918_ clknet_leaf_101_wb_clk_i _03468_ _01738_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_94_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08164__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1180 net1182 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__buf_4
Xfanout1191 net1194 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_2
XFILLER_0_20_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08651_ net1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\] net925
+ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__and3_1
XANTENNA__09900__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17849_ clknet_leaf_106_wb_clk_i net2851 _01669_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17832__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08582_ _04835_ _04837_ _04839_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09113__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12365__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10274__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13748__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09203_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] net909
+ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09134_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] net887
+ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18017__1594 vssd1 vssd1 vccd1 vccd1 net1594 _18017__1594/LO sky130_fd_sc_hd__conb_1
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12971__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\] net867
+ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14182__C _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14173__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold630 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold663 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\] vssd1 vssd1 vccd1 vccd1
+ net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout861_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] net898 vssd1
+ vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__and3_1
X_18186__1560 vssd1 vssd1 vccd1 vccd1 _18186__1560/HI net1560 sky130_fd_sc_hd__conb_1
X_08918_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\] net898
+ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__and3_1
XANTENNA__12203__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] net654 net623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__a22o_1
Xhold1330 _03450_ vssd1 vssd1 vccd1 vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08155__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1341 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1352 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2968 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1363 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] vssd1 vssd1 vccd1 vccd1
+ net2979 sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\] net850 vssd1
+ vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__and3_1
XANTENNA__13245__D net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net2990
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 team_01_WB.instance_to_wrap.cpu.K0.code\[3\] vssd1 vssd1 vccd1 vccd1 net3012
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11860_ _07850_ _07976_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__or2_1
XANTENNA__08917__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__B1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10811_ net543 _07074_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__and2_1
X_11791_ net2132 net284 net479 vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13530_ net1066 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _03879_ _03880_
+ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10742_ _05583_ _05515_ net502 vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10673_ _06778_ _06936_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nor2_1
X_13461_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _05550_ vssd1 vssd1
+ vccd1 vccd1 _03814_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15200_ net1273 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
X_12412_ net2596 net219 net420 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
XANTENNA__09748__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16180_ clknet_leaf_91_wb_clk_i _01848_ _00048_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_13392_ net2858 net329 net353 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1
+ vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08652__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15131_ net1300 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12343_ net2953 net225 net492 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__mux2_1
XANTENNA__08630__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15062_ net1303 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
X_12274_ net2308 net288 net431 vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14013_ team_01_WB.EN_VAL_REG net2927 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11225_ _07487_ _07488_ _05891_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__o21ba_1
X_18070__1444 vssd1 vssd1 vccd1 vccd1 _18070__1444/HI net1444 sky130_fd_sc_hd__conb_1
XANTENNA__10125__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ _07339_ _07419_ net535 vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__mux2_1
XANTENNA__17855__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] net621 net617 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11518__A team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15964_ net1336 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__inv_2
X_11087_ _06178_ _07350_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12113__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17703_ clknet_leaf_72_wb_clk_i _03263_ _01542_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08146__B2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[4\] net844 vssd1
+ vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__and3_1
X_14915_ net1220 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15895_ net1350 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11952__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17634_ clknet_leaf_143_wb_clk_i _03194_ _01497_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14846_ net1384 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09422__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17565_ clknet_leaf_127_wb_clk_i _03125_ _01428_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14777_ net1337 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XANTENNA__08449__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ net2000 net268 net468 vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16516_ clknet_leaf_75_wb_clk_i _02144_ _00379_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13728_ _04464_ _04025_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ clknet_leaf_26_wb_clk_i _03056_ _01359_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16447_ clknet_leaf_77_wb_clk_i net2184 _00310_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12783__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13659_ net773 _07368_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10008__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16378_ clknet_leaf_110_wb_clk_i net1809 _00246_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12953__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18117_ net1491 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15329_ net1291 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11700__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08621__A2 _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14155__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ net1610 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_111_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09096__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10035__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 _03563_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_4
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_6
XANTENNA__09582__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09393__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\] net858 vssd1
+ vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__and3_1
Xfanout428 _08024_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13627__B _07551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 _08021_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_6
XANTENNA__09824__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] net651 _06000_
+ _06001_ _06009_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12023__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08703_ net971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] net929 vssd1
+ vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__and3_1
X_09683_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] net874
+ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__and3_1
XANTENNA__08688__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout275_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18010__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08634_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] net665 net641 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08565_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\] net658 net609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout442_A _08021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1184_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__A2_N net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08496_ net1106 net1108 net1111 net1114 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_71_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12693__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16602__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08860__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09568__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12944__B2 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] net879
+ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08612__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] net897
+ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16752__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold460 _02080_ vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net330 _07070_ _07096_ net521 net532 vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__a221o_1
Xhold493 team_01_WB.instance_to_wrap.a1.ADR_I\[20\] vssd1 vssd1 vccd1 vccd1 net2109
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09734__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout940 net941 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_8
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_2
Xfanout962 net964 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
Xfanout973 net976 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net1009 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlymetal6s2s_1
X_12961_ net1670 net604 net586 _03647_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08679__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 _02130_ vssd1 vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] vssd1 vssd1 vccd1 vccd1
+ net2787 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ net1373 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net2110 net282 net475 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
X_15680_ net1273 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
Xhold1193 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] net1056 net366 _03597_
+ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a22o_1
XANTENNA__08647__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17258__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ net1371 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _07851_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11435__A1 _04592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17350_ clknet_leaf_141_wb_clk_i _02910_ _01213_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ net1331 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ net2515 net200 net479 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16301_ clknet_leaf_112_wb_clk_i _01935_ _00169_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13513_ _03755_ _03865_ _03756_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a21bo_1
X_17281_ clknet_leaf_137_wb_clk_i _02841_ _01144_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10725_ _06978_ _06987_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__or2_2
XFILLER_0_82_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14493_ net1358 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XANTENNA__16282__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16232_ clknet_leaf_37_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[13\]
+ _00100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13444_ _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10656_ _05485_ _06919_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__nand2_1
XANTENNA__08813__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16163_ clknet_leaf_90_wb_clk_i _01831_ _00031_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13375_ net2341 net328 net352 net1062 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
XANTENNA__12108__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08603__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] _04716_ _06850_ vssd1 vssd1
+ vccd1 vccd1 _06851_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11012__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15114_ net1223 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
X_12326_ net3134 net261 net429 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16094_ net1371 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11947__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ net1225 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12257_ net2488 net315 net437 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__mux2_1
XANTENNA__10851__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13360__A1 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ net520 _07210_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__nand2_2
X_12188_ net2078 net267 net445 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13447__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ _06141_ _06211_ net506 vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__mux2_1
X_16996_ clknet_leaf_128_wb_clk_i _02556_ _00859_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13112__A1 _06559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15947_ net1396 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12778__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ net1393 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17617_ clknet_leaf_20_wb_clk_i _03177_ _01480_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14829_ net1347 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] net1626 net1047 vssd1 vssd1
+ vccd1 vccd1 _03397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17548_ clknet_leaf_45_wb_clk_i _03108_ _01411_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08281_ net2138 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17479_ clknet_leaf_130_wb_clk_i _03039_ _01342_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11711__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09819__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12018__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14128__B1 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11857__S net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout203 _07888_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_1
Xfanout214 _08007_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13351__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 _07915_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout236 net237 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout247 net249 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
X_09804_ _06048_ _06056_ _06057_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or4_1
XANTENNA__10062__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout269 _07962_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09851__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\] net843 vssd1
+ vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17400__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12688__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout657_A _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09666_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] net848
+ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__and3_1
XANTENNA__11665__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ net713 _04873_ _04877_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__or4_2
X_09597_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\] net891 vssd1
+ vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout824_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17550__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08548_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] net731 net695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ net1084 net886 vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__and2_2
XFILLER_0_33_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09298__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ _06772_ _06773_ net578 vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__mux2_1
X_11490_ team_01_WB.instance_to_wrap.cpu.DM0.dhit _07724_ vssd1 vssd1 vccd1 vccd1
+ _07739_ sky130_fd_sc_hd__and2_2
XFILLER_0_11_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10441_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] net628 net618 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\]
+ _06704_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__a221o_1
XANTENNA__10237__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09794__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ net2501 net2441 net826 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
X_10372_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] net747 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13590__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ net2583 net228 net451 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__mux2_1
XANTENNA__10943__A3 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ net356 _03713_ _03714_ net836 net1700 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09546__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net3070 net287 net459 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold290 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09010__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16850_ clknet_leaf_22_wb_clk_i _02410_ _00713_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15801_ net1191 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
Xfanout770 _04626_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_4
Xfanout781 _04622_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_2
X_16781_ clknet_leaf_20_wb_clk_i _02341_ _00644_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13993_ _04160_ _03554_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12598__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15732_ net1237 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ net1899 net604 net586 _03635_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11656__B2 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08377__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08808__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15663_ net1246 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
X_12875_ net2275 net607 _03584_ net589 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
X_17402_ clknet_leaf_36_wb_clk_i _02962_ _01265_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14614_ net1378 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11826_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07853_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09077__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15594_ net1202 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16798__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17333_ clknet_leaf_9_wb_clk_i _02893_ _01196_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14545_ net1319 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11757_ net774 _07890_ _07892_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__o21ai_4
XANTENNA__08824__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13222__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17264_ clknet_leaf_23_wb_clk_i _02824_ _01127_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ net544 _06970_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__nand2_1
X_14476_ net1335 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
X_11688_ net2816 _07837_ net36 vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a21o_1
XANTENNA__09639__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18165__1539 vssd1 vssd1 vccd1 vccd1 _18165__1539/HI net1539 sky130_fd_sc_hd__conb_1
XFILLER_0_71_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16215_ clknet_leaf_117_wb_clk_i _01882_ _00083_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__08543__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] _06348_ vssd1 vssd1 vccd1
+ vccd1 _03780_ sky130_fd_sc_hd__nand2_1
XANTENNA__15938__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17195_ clknet_leaf_60_wb_clk_i _02755_ _01058_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10639_ _05963_ _06030_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13581__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16146_ net1321 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09936__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13358_ net29 net802 _03747_ net2808 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
XANTENNA__08840__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ net2879 net228 net427 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
X_16077_ net1347 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__inv_2
X_13289_ net97 net812 net598 net1885 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16178__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15028_ net1241 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17423__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09671__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13097__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13905__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16979_ clknet_leaf_49_wb_clk_i _02539_ _00842_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
XFILLER_0_36_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09520_ _05780_ _05781_ _05782_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__or4_1
XANTENNA__12301__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09390__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09451_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] net731 net711 _05713_
+ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08402_ net1152 net1154 net1148 net1150 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__and4bb_4
X_09382_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\] net742 net705 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12072__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08333_ net2626 net2710 net1044 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XANTENNA__10756__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__mux2_1
XANTENNA__10622__A2 _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11262__A1_N _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08195_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] _04592_ _04567_ vssd1 vssd1 vccd1
+ vccd1 _04595_ sky130_fd_sc_hd__mux2_1
XANTENNA__10057__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08750__A _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1314_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 _04484_ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11335__B1 _07598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13875__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11886__A1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13088__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] net689 _05967_
+ _05972_ _05977_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11638__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10520__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10990_ _05417_ net342 net335 _05416_ net333 vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16940__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[11\] net696 _05895_
+ _05903_ _05906_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12660_ net2031 net294 net394 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11611_ net497 _07820_ net2163 net838 vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ net2361 net260 net401 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__mux2_1
XANTENNA__13260__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14330_ net3138 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _07706_ _07739_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09459__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\] _04244_ _04249_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\]
+ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__a221o_1
X_11473_ _04463_ _07725_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ net1359 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__inv_2
XANTENNA_input70_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net2840 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\] net819 vssd1 vssd1
+ vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10424_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\] net715 net700 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16320__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14192_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\] _04246_ _04346_ _04348_
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__17446__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13143_ net2455 net1767 net831 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10355_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\] net927
+ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10286_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\] _04754_
+ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__and3_1
X_13074_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\] _03702_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__mux2_1
X_17951_ clknet_leaf_108_wb_clk_i _03501_ _01771_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09194__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12025_ net2060 net315 net464 vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
X_16902_ clknet_leaf_139_wb_clk_i _02462_ _00765_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12332__D team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17882_ clknet_leaf_78_wb_clk_i _03432_ _01702_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09491__A _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16833_ clknet_leaf_135_wb_clk_i _02393_ _00696_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09922__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14276__C1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12121__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ clknet_leaf_10_wb_clk_i _02324_ _00627_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13976_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\]
+ net584 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15715_ net1222 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__08538__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ net1026 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\] vssd1 vssd1 vccd1
+ vccd1 _03623_ sky130_fd_sc_hd__or2_1
X_16695_ clknet_leaf_11_wb_clk_i _02255_ _00558_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11960__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15646_ net1316 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12858_ net2108 net294 net369 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10584__C_N team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07855_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\]
+ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15577_ net1190 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
X_12789_ net1933 net259 net377 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17316_ clknet_leaf_128_wb_clk_i _02876_ _01179_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14528_ net1322 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XANTENNA__11801__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09369__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17247_ clknet_leaf_1_wb_clk_i _02807_ _01110_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14459_ net1390 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XANTENNA__12791__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10308__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17178_ clknet_leaf_34_wb_clk_i _02738_ _01041_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11565__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16129_ net1397 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16813__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13306__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08951_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] net950
+ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_122_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08882_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\] net925
+ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16963__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12031__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09503_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] net948 vssd1
+ vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11096__A2 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09434_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] net920 vssd1
+ vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09365_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] net917
+ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout522_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1264_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08316_ net3120 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\] net1039 vssd1 vssd1
+ vccd1 vccd1 _03431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[14\] net937
+ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09749__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _04554_ _04565_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09213__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout891_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16493__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12206__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10140_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\] _04641_ net719 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\]
+ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__13248__D net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
X_10071_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\] net751 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11859__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09742__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18164__1538 vssd1 vssd1 vccd1 vccd1 _18164__1538/HI net1538 sky130_fd_sc_hd__conb_1
X_13830_ team_01_WB.instance_to_wrap.cpu.c0.count\[14\] team_01_WB.instance_to_wrap.cpu.c0.count\[13\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[12\] team_01_WB.instance_to_wrap.cpu.c0.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__or4b_1
XFILLER_0_98_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13761_ net1672 _04071_ net783 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__mux2_1
XANTENNA__11784__A1_N net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__S net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ net539 _07133_ _07234_ _06996_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__a211o_1
XANTENNA__11780__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15500_ net1265 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
X_12712_ net3108 net278 net383 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16480_ clknet_leaf_109_wb_clk_i _02108_ _00343_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\]
+ sky130_fd_sc_hd__dfstp_1
X_13692_ _07710_ _07774_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ net1182 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
X_12643_ net2898 net221 net392 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18150_ net1524 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
XFILLER_0_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15362_ net1311 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12574_ net2428 net227 net399 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__mux2_1
XANTENNA__09189__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17101_ clknet_leaf_21_wb_clk_i _02661_ _00964_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11795__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14313_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] _04450_ net1991 vssd1
+ vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ net1063 _07762_ _07763_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18081_ net1455 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15293_ net1280 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
XANTENNA__08660__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16836__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ clknet_leaf_45_wb_clk_i _02592_ _00895_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10128__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\] _04249_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a221o_1
X_11456_ _07708_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__inv_2
XANTENNA__08390__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10407_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] net920 vssd1
+ vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] _04261_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a221o_1
XANTENNA__12116__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__A2 _06995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ net533 _07258_ _07650_ net321 vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ net821 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
X_10338_ _06180_ _06599_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10770__A1 _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13736__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13057_ _05133_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__o21a_1
X_17934_ clknet_leaf_101_wb_clk_i _03484_ _01754_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\]
+ sky130_fd_sc_hd__dfstp_1
X_10269_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\] net888 vssd1
+ vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__and3_1
Xfanout1340 net1349 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__buf_4
X_12008_ net2285 net231 net464 vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1351 net1360 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__buf_4
Xfanout1362 net1365 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__clkbuf_4
X_17865_ clknet_leaf_108_wb_clk_i _03415_ _01685_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1373 net1379 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__buf_4
Xfanout1384 net1385 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__buf_4
Xfanout1395 net1398 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__buf_4
XFILLER_0_89_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16816_ clknet_leaf_23_wb_clk_i _02376_ _00679_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17796_ clknet_leaf_70_wb_clk_i _03353_ _01617_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13959_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__or4b_1
X_16747_ clknet_leaf_51_wb_clk_i _02307_ _00610_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12786__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16678_ clknet_leaf_87_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_dhit _00541_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.dhit sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09691__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11703__B _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15629_ net1217 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09150_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] net668 _05409_ _05413_
+ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10589__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08101_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] _04495_ team_01_WB.instance_to_wrap.cpu.f0.num\[9\]
+ _04476_ _04517_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09081_ _05310_ _05344_ net583 vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10038__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 _04463_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput50 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput61 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput72 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
Xhold801 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09827__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold812 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold834 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12026__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold856 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10210__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold867 _03490_ vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold878 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09983_ _06211_ _06245_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__nand2_1
Xhold889 _03423_ vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ _05187_ _05188_ _05189_ _05190_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout1012_A _04484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1501 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] vssd1 vssd1 vccd1 vccd1
+ net3128 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09562__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] net660 _05115_ _05116_
+ _05122_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a2111o_1
Xhold1523 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net3139 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout472_A _08010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1534 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15861__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1556 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3183 sky130_fd_sc_hd__dlygate4sd3_1
X_08796_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] net648 net633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
Xhold1578 team_01_WB.instance_to_wrap.cpu.f0.num\[1\] vssd1 vssd1 vccd1 vccd1 net3194
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1381_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08475__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17291__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08906__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] net655 net622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a22o_1
XANTENNA__08890__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout904_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16859__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13766__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09348_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] net638 _05591_ _05596_
+ _05606_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11777__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\] net661 _05520_ _05528_
+ _05530_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11241__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15101__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ net537 _07472_ _07573_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ net2743 net316 net431 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09737__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ _06029_ net337 net331 _06028_ _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11172_ net511 _07015_ _07017_ _07435_ net524 vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__o311a_1
XANTENNA__10752__A1 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16239__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10123_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] net963 vssd1
+ vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__and3_1
X_15980_ net1385 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10054_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__inv_2
X_14931_ net1186 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17650_ clknet_leaf_40_wb_clk_i _03210_ _01513_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14862_ net1346 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16389__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14246__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10411__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13813_ net2025 _04511_ _04559_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1
+ vccd1 vccd1 _01829_ sky130_fd_sc_hd__a22o_1
X_16601_ clknet_leaf_104_wb_clk_i _02229_ _00464_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_17581_ clknet_leaf_19_wb_clk_i _03141_ _01444_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14793_ net1333 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16532_ clknet_leaf_56_wb_clk_i _02160_ _00395_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ _07720_ _07752_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10956_ _05621_ _06036_ _07205_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08385__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08816__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16463_ clknet_leaf_76_wb_clk_i net1772 _00326_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13675_ net770 _03999_ net969 vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10887_ _07136_ _07141_ _07150_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11015__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18202_ net1576 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17784__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15414_ net1305 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ net2248 net308 net398 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16394_ clknet_leaf_102_wb_clk_i _02022_ _00257_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18133_ net1507 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
XFILLER_0_108_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15345_ net1200 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
X_12557_ net1855 net300 net405 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13230__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11508_ _04467_ _07719_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__nand2_1
XANTENNA__10440__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18064_ net1438 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12980__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15276_ net1252 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12488_ net2350 net305 net412 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold108 _01955_ vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17015_ clknet_leaf_12_wb_clk_i _02575_ _00878_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 _01997_ vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\] _04264_ _04276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\]
+ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a221o_1
XANTENNA__15946__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11439_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ _04598_ _07683_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14158_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\] _04252_ _04315_ _04317_
+ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13109_ net2156 net837 net357 _03724_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a22o_1
XANTENNA__17164__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14089_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\] _04249_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\]
+ _04248_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17917_ clknet_leaf_104_wb_clk_i _03467_ _01737_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_59_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15681__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1170 net1172 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
X_08650_ net1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] net927
+ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__and3_1
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_4
Xfanout1192 net1194 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_4
X_17848_ clknet_leaf_98_wb_clk_i net1867 _01668_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] net662 _04829_
+ _04842_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17779_ clknet_leaf_116_wb_clk_i _03337_ _01600_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11714__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13996__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] net904
+ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13748__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11759__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ net1075 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] net870
+ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__and3_1
XANTENNA__08624__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09064_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] net842
+ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and3_1
XANTENNA__12971__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18163__1537 vssd1 vssd1 vccd1 vccd1 _18163__1537/HI net1537 sky130_fd_sc_hd__conb_1
XANTENNA__08234__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08461__C _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14182__D _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10065__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold642 net130 vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1227_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\] vssd1 vssd1 vccd1 vccd1
+ net2269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09854__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold664 _02034_ vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09966_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] net873 vssd1
+ vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08917_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\] net879
+ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__and3_1
XANTENNA__09292__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] net869 vssd1
+ vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1320 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\] vssd1 vssd1 vccd1 vccd1
+ net2936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1331 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] vssd1 vssd1 vccd1 vccd1
+ net2947 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10498__B1 _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1342 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2958 sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] net898
+ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__and3_1
Xhold1353 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2969 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1364 _02089_ vssd1 vssd1 vccd1 vccd1 net2980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14228__A2 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1375 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2991 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10231__C net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1386 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\] vssd1 vssd1 vccd1 vccd1
+ net3002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1397 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08779_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] net762 _05041_ _05042_
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a22o_4
XANTENNA__09104__A1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ net549 net538 vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11790_ net775 _07917_ _07918_ _07919_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__09655__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _05718_ net548 net503 vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ _03793_ _03810_ _03812_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o21ai_1
X_10672_ _06828_ _06807_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__nand2b_1
XANTENNA__17037__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ net2187 net282 net419 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13391_ net2796 net327 net351 net1065 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XANTENNA__08615__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15130_ net1305 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12342_ net3026 net227 net490 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09467__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ net1173 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12273_ net2141 net232 net433 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
X_14012_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\] _04192_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.lcd_en sky130_fd_sc_hd__a21oi_1
XANTENNA__10406__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09764__A _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _05823_ net343 net336 _05822_ net333 vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__a221o_1
XANTENNA__09040__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11155_ _07108_ _07113_ net529 vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__mux2_1
XANTENNA__10703__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10106_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\] net659 _06355_ _06364_
+ _06367_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12478__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15963_ net1337 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__inv_2
X_11086_ _06141_ _06175_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13675__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17702_ clknet_leaf_72_wb_clk_i _03262_ _01541_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10037_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\] net884 vssd1
+ vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__and3_1
X_14914_ net1290 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
X_15894_ net1356 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__A1 _06870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14219__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ clknet_leaf_136_wb_clk_i _03193_ _01496_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09930__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14845_ net1359 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11534__A team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15006__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14776_ net1333 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17564_ clknet_leaf_13_wb_clk_i _03124_ _01427_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11988_ net2393 net272 net467 vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_1
XANTENNA__13928__A_N net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09646__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08546__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ _04558_ _04020_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__or3_1
X_16515_ clknet_leaf_101_wb_clk_i net2035 _00378_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _06033_ _06604_ _05761_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__a21o_1
X_17495_ clknet_leaf_12_wb_clk_i _03055_ _01358_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16446_ clknet_leaf_80_wb_clk_i _02074_ _00309_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_13658_ _07977_ _03986_ net188 vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08843__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ net2311 net285 net396 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
X_16377_ clknet_leaf_111_wb_clk_i net1774 _00245_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13589_ net773 _07625_ net966 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15328_ net1276 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
X_18116_ net1490 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_26_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12953__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_134_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15259_ net1316 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
X_18047_ net1609 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09674__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09031__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09820_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] net898 vssd1
+ vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__and3_1
Xfanout407 _03562_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_8
Xfanout418 _08029_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11709__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12304__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 _08024_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_8
X_09751_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] net639 net609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__a22o_1
XANTENNA__13666__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12332__A_N _07834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] net917
+ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__and3_1
X_09682_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\] net866
+ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08633_ _04890_ _04892_ _04894_ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13418__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] net759 _04826_ _04827_
+ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a22o_2
XFILLER_0_72_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08495_ net1072 net870 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout435_A _08022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09849__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08753__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] net576 net577 vssd1 vssd1
+ vccd1 vccd1 _05380_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12944__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09047_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\] net886
+ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10226__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold461 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold472 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold483 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12214__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold494 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10523__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10183__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout930 net934 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_4
Xfanout941 _04657_ vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_6
X_09949_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] net667 vssd1 vssd1
+ vccd1 vccd1 _06213_ sky130_fd_sc_hd__or2_2
Xfanout952 _04644_ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_6
Xfanout963 _04638_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_4
Xfanout974 net976 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 net992 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
X_12960_ _03582_ _03645_ _03646_ team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net1009 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11132__A1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1150 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1161 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ net3182 net223 net477 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 _03485_ vssd1 vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] _07153_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03597_ sky130_fd_sc_hd__mux2_1
Xhold1183 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\] vssd1 vssd1 vccd1 vccd1
+ net2810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ net1375 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ net1976 net266 net481 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ net1331 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ net777 _07903_ _07904_ _07905_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13512_ _03757_ _03758_ _03862_ _04955_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a32o_1
X_16300_ clknet_leaf_112_wb_clk_i _01934_ _00168_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17280_ clknet_leaf_2_wb_clk_i _02840_ _01143_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ _06978_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__nor2_1
X_14492_ net1361 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16231_ clknet_leaf_37_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[12\]
+ _00099_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[12\] sky130_fd_sc_hd__dfrtp_1
X_13443_ _05924_ _03794_ _03795_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_125_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10655_ _06899_ _06904_ _06918_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__a21o_2
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08382__B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16162_ clknet_leaf_90_wb_clk_i _01830_ _00030_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13374_ net2533 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1
+ vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XANTENNA__16577__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09197__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10586_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] _04628_ _04633_ vssd1 vssd1
+ vccd1 vccd1 _06850_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09800__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15113_ net1221 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
X_12325_ net2729 net299 net430 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
X_16093_ net1348 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__inv_2
XANTENNA__12913__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15044_ net1270 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XANTENNA__09494__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ net2516 net303 net437 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ net537 _07470_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12124__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ net2937 net270 net443 vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__mux2_1
XANTENNA__17972__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ net331 _07400_ _07401_ _06246_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__a31o_1
XANTENNA__11248__B _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__B _06415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16995_ clknet_leaf_132_wb_clk_i _02555_ _00858_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11963__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15946_ net1396 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _06991_ _07074_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A1 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09867__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17202__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18162__1536 vssd1 vssd1 vccd1 vccd1 _18162__1536/HI net1536 sky130_fd_sc_hd__conb_1
X_15877_ net1392 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17616_ clknet_leaf_30_wb_clk_i _03176_ _01479_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10882__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14828_ net1341 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12794__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17547_ clknet_leaf_51_wb_clk_i _03107_ _01410_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08827__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14759_ net1221 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17352__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09669__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17478_ clknet_leaf_140_wb_clk_i _03038_ _01341_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16429_ clknet_leaf_78_wb_clk_i _02057_ _00292_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11711__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13351__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout204 _07888_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
Xfanout215 _07943_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
Xfanout226 _07911_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
XFILLER_0_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout237 _07893_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
X_09803_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] _04646_ net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__a22o_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_2
Xfanout259 _07989_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
XANTENNA_fanout385_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net1008 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] net881 vssd1
+ vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09665_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\] net880
+ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout552_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09570__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1294_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ _04867_ _04868_ _04878_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09596_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] net863 vssd1
+ vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08547_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\] net944 vssd1
+ vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08818__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13811__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ net1107 net1112 net1114 net1109 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_114_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17845__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08914__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12209__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10518__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10440_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\] net640 net638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09243__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11050__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] net750 net703 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\]
+ _06623_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ net2173 net201 net451 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13090_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\] net1026 vssd1 vssd1 vccd1
+ vccd1 _03714_ sky130_fd_sc_hd__or2_1
XANTENNA__09745__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13342__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ net3220 net230 net460 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold280 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18109__1483 vssd1 vssd1 vccd1 vccd1 _18109__1483/HI net1483 sky130_fd_sc_hd__conb_1
XANTENNA__17225__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout760 net761 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
X_15800_ net1242 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__inv_2
Xfanout771 net773 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_2
Xfanout782 net784 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
X_16780_ clknet_leaf_47_wb_clk_i _02340_ _00643_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13992_ net1403 _04160_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout793 _04223_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12943_ net364 _03633_ _03634_ net1053 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a32o_1
X_15731_ net1189 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08377__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08521__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15662_ net1230 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_12874_ net1055 team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] net606 vssd1 vssd1
+ vccd1 vccd1 _03585_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17401_ clknet_leaf_125_wb_clk_i _02961_ _01264_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11825_ net2118 net277 net480 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14613_ net1375 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
X_15593_ net1210 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XANTENNA__12908__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14544_ net1322 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17332_ clknet_leaf_7_wb_clk_i _02892_ _01195_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11756_ net675 _07152_ _07891_ net781 vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ net542 net531 _06953_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__and3_4
X_14475_ net1335 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17263_ clknet_leaf_18_wb_clk_i _02823_ _01126_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11687_ net2646 net1169 net37 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a21o_1
XANTENNA__12119__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13426_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _06278_ vssd1 vssd1 vccd1
+ vccd1 _03779_ sky130_fd_sc_hd__and2_1
X_16214_ clknet_leaf_117_wb_clk_i _01881_ _00082_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ sky130_fd_sc_hd__dfstp_2
X_17194_ clknet_leaf_41_wb_clk_i _02754_ _01057_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13030__A1 _04902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10638_ _05758_ _05760_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ net1321 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__inv_2
XANTENNA__11958__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ net30 net800 net595 net2320 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__o22a_1
XANTENNA__13581__A2 _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap916 _04677_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_2
X_10569_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10395__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ net2102 net198 net427 vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
X_16076_ net1403 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__inv_2
X_13288_ net100 net812 net597 net1832 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08332__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15027_ net1189 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13333__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ net3206 net235 net435 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10163__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10147__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__A1 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12789__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13474__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13097__A1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17718__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16978_ clknet_leaf_22_wb_clk_i _02538_ _00841_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15929_ net1351 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09450_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\] net753 _05690_
+ _05698_ _05700_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_56_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16742__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\] net931
+ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and3_1
XANTENNA__17868__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09381_ _05641_ _05642_ _05643_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11722__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ net2504 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\] net1038 vssd1 vssd1
+ vccd1 vccd1 _03415_ sky130_fd_sc_hd__mux2_1
XANTENNA__09399__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10083__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux2_1
XANTENNA__12029__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__A3 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08194_ _04568_ _04593_ _04594_ net553 net1667 vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__a32o_1
XANTENNA__13021__A1 _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08579__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16025__A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10386__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17248__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18036__1602 vssd1 vssd1 vccd1 vccd1 net1602 _18036__1602/LO sky130_fd_sc_hd__conb_1
XFILLER_0_125_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13324__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1307_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11889__A2_N net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12699__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16272__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17398__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13088__A1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\] net716 _05965_ _05973_
+ _05974_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08909__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09648_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\] net688 _05894_
+ _05897_ _05898_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09579_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\] net729 net706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11610_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[21\] net572 vssd1 vssd1 vccd1
+ vccd1 _07820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15104__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12590_ net3192 net298 net402 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08644__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net1065 _07706_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13548__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\] _04272_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__a22o_1
X_11472_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] team_01_WB.instance_to_wrap.cpu.f0.i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08941__A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13211_ net2660 net2617 net825 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
X_10423_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\] net748 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\]
+ _06678_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__a221o_1
X_14191_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\] _04239_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\]
+ _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18161__1535 vssd1 vssd1 vccd1 vccd1 _18161__1535/HI net1535 sky130_fd_sc_hd__conb_1
XFILLER_0_81_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13142_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
XANTENNA_input63_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\] net925 vssd1
+ vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13073_ _05549_ net570 net359 vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o21a_1
X_17950_ clknet_leaf_101_wb_clk_i _03500_ _01770_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__16615__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10285_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] _04749_ net615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\]
+ _06548_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10414__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ net2151 net304 net464 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
X_16901_ clknet_leaf_132_wb_clk_i _02461_ _00764_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09772__A _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17881_ clknet_leaf_109_wb_clk_i _03431_ _01701_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08742__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_137_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16832_ clknet_leaf_140_wb_clk_i _02392_ _00695_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13079__A1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12402__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14276__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _04849_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_2
XANTENNA__16765__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16763_ clknet_leaf_37_wb_clk_i _02323_ _00626_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11629__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] _04153_ _04165_ net1170
+ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__o211a_2
XFILLER_0_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15714_ net1313 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
X_12926_ net1026 _07520_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nand2_1
X_16694_ clknet_leaf_31_wb_clk_i _02254_ _00557_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ net1282 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12857_ net2119 net307 net369 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11808_ net1920 net252 net481 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ net2002 net298 net378 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
X_15576_ net1242 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17315_ clknet_leaf_132_wb_clk_i _02875_ _01178_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11262__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11261__B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14527_ net1314 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
X_11739_ net674 _07600_ _07877_ net781 vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10158__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09207__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17246_ clknet_leaf_139_wb_clk_i _02806_ _01109_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14458_ net1390 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
XANTENNA__14200__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _06717_ vssd1 vssd1
+ vccd1 vccd1 _03762_ sky130_fd_sc_hd__nor2_1
X_14389_ net1327 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17177_ clknet_leaf_16_wb_clk_i _02737_ _01040_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10368__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16128_ net1395 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16295__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] net957
+ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__and3_1
XANTENNA__13306__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15684__A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16059_ net1413 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09682__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13916__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08881_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\] net941
+ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08194__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08733__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14267__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10540__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12817__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09502_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\] net943 vssd1
+ vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11096__A3 _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\] net953 vssd1
+ vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout250_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] net924
+ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__and3_1
XANTENNA__13242__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08315_ net3052 net3212 net1049 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18108__1482 vssd1 vssd1 vccd1 vccd1 _18108__1482/HI net1482 sky130_fd_sc_hd__conb_1
X_09295_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\] net926
+ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout515_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1257_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09857__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08246_ net3175 net3002 net1039 vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13545__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ net1803 net553 _04568_ _04578_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a22o_1
XANTENNA__16638__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09295__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08972__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XANTENNA__11308__A1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10234__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__09592__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[3\] net750 _04656_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08724__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12222__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10531__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13760_ net484 _07717_ _04068_ _04070_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__a31o_1
X_10972_ _05348_ net340 net338 _05347_ _07235_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__o221a_1
XANTENNA__08936__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12711_ net2992 net253 net385 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__mux2_1
X_13691_ _03744_ _04012_ _04013_ net1166 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15430_ net1278 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
X_12642_ net1942 net282 net391 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ net1290 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12573_ net2845 net198 net399 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17100_ clknet_leaf_44_wb_clk_i _02660_ _00963_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11524_ net1063 _07732_ _07761_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14312_ net2933 _04450_ _04452_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o21a_1
XANTENNA__10409__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15292_ net1232 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
X_18080_ net1454 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_110_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17031_ clknet_leaf_130_wb_clk_i _02591_ _00894_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14243_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] _04244_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\]
+ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a22o_1
X_11455_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] team_01_WB.instance_to_wrap.cpu.f0.i\[13\]
+ _07706_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17563__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11547__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10706__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10406_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\] net961
+ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__and3_1
X_14174_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\] _04258_ _04278_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\]
+ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11386_ net525 _07187_ _07649_ net537 vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ net823 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
XANTENNA__08963__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ _06319_ _06597_ _06600_ _06599_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13056_ net1877 net834 net355 _03690_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
X_17933_ clknet_leaf_105_wb_clk_i _03483_ _01753_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\]
+ sky130_fd_sc_hd__dfstp_1
X_10268_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] net873 vssd1
+ vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09933__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__B1 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1330 net1337 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__buf_4
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ net3186 net237 net463 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__mux2_1
XANTENNA__08715__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1341 net1342 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__buf_4
XANTENNA__12132__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1352 net1360 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__buf_4
X_17864_ clknet_leaf_99_wb_clk_i _03414_ _01684_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10199_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] net926 vssd1
+ vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__and3_1
XANTENNA__14249__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1363 net1364 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1374 net1379 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__clkbuf_4
X_16815_ clknet_leaf_18_wb_clk_i _02375_ _00678_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1385 net1388 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__buf_4
Xfanout1396 net1398 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__buf_4
X_17795_ clknet_leaf_70_wb_clk_i _03352_ _01616_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11971__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16746_ clknet_leaf_42_wb_clk_i _02306_ _00609_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13958_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__or4b_1
XANTENNA__08846__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09140__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\] vssd1 vssd1 vccd1
+ vccd1 _03610_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16677_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[31\]
+ _00540_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13889_ net2252 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[2\]
+ sky130_fd_sc_hd__and2_1
X_18035__1601 vssd1 vssd1 vccd1 vccd1 net1601 _18035__1601/LO sky130_fd_sc_hd__conb_1
XFILLER_0_134_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15628_ net1265 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17093__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11703__C _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ net1180 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08100_ _04464_ team_01_WB.instance_to_wrap.cpu.f0.num\[25\] team_01_WB.instance_to_wrap.cpu.f0.num\[1\]
+ _04482_ _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a221o_1
XANTENNA__12983__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17906__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09080_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] net666 _05340_ _05343_
+ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__o22a_4
XFILLER_0_12_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08031_ net1061 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__inv_2
Xinput40 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
X_17229_ clknet_leaf_50_wb_clk_i _02789_ _01092_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12307__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput62 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
Xhold802 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold813 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold824 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold835 team_01_WB.instance_to_wrap.cpu.f0.num\[29\] vssd1 vssd1 vccd1 vccd1 net2451
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09982_ _06211_ _06245_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nor2_1
Xhold868 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold879 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08933_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\] net643 _05196_
+ net672 vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__B1 _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1502 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12042__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] _04755_ _05101_
+ _05114_ net672 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a2111o_1
Xhold1513 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\] vssd1 vssd1 vccd1 vccd1
+ net3129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1005_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1524 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1 vccd1
+ net3151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08459__C net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1546 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3173 sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] net655 net629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1568 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11881__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1579 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18160__1534 vssd1 vssd1 vccd1 vccd1 _18160__1534/HI net1534 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1374_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _05676_ _05677_ _05678_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__nor4_1
XFILLER_0_133_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09347_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\] net630 _05587_
+ _05590_ _05595_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17586__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10229__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] net637 _05532_
+ _05534_ _05537_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_118_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08491__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08922__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ net1713 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10526__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ _06027_ net335 vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__nand2_1
XANTENNA__14191__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11171_ net511 _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10122_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] net744 net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a22o_1
XANTENNA__09355__C1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ _06277_ net547 vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nor2_1
X_14930_ net1188 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XANTENNA__10504__A2 _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1346 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11791__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16600_ clknet_leaf_66_wb_clk_i _02228_ _00463_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13812_ net1747 net784 _07681_ _04109_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__o22a_1
X_17580_ clknet_leaf_46_wb_clk_i _03140_ _01443_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14792_ net1327 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
X_16531_ clknet_leaf_61_wb_clk_i _02159_ _00394_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13743_ _04555_ _04056_ team_01_WB.instance_to_wrap.cpu.f0.next_write_i vssd1 vssd1
+ vccd1 vccd1 _04057_ sky130_fd_sc_hd__o21a_1
X_10955_ _06036_ _07202_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17929__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16462_ clknet_leaf_86_wb_clk_i _02090_ _00325_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13674_ net770 _07426_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10886_ net545 _07145_ _07148_ _07149_ _07147_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18201_ net1575 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
X_15413_ net1175 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
X_12625_ net2819 net313 net397 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XANTENNA__15499__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16393_ clknet_leaf_73_wb_clk_i _02021_ _00256_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_38_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ net1506 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
XANTENNA__12965__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15344_ net1262 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ net2823 net242 net405 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11507_ net1062 _07750_ _07751_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18063_ net1437 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
X_12487_ net1932 net264 net412 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XANTENNA__12127__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ net1207 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold109 net112 vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17014_ clknet_leaf_33_wb_clk_i _02574_ _00877_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10991__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11438_ _07694_ net1649 _07685_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14226_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\] _04275_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13747__A team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_104_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14157_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[98\] _04250_ _04276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\]
+ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a221o_1
XANTENNA__17309__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ net510 _07055_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13108_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] _06450_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14088_ _04226_ net788 _04241_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__and3_4
XANTENNA__08340__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__C net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17916_ clknet_leaf_81_wb_clk_i _03466_ _01736_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_13039_ _06716_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__o21a_1
XANTENNA__10171__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18107__1481 vssd1 vssd1 vccd1 vccd1 _18107__1481/HI net1481 sky130_fd_sc_hd__conb_1
Xfanout1160 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1160
+ sky130_fd_sc_hd__buf_2
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17459__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09960__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17847_ clknet_leaf_86_wb_clk_i _03397_ _01667_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout1182 net1185 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_4
XANTENNA__12797__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_2
XFILLER_0_55_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] net646 net638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\]
+ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__a221o_1
X_17778_ clknet_leaf_116_wb_clk_i _03336_ _01599_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10259__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09113__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16729_ clknet_leaf_16_wb_clk_i _02289_ _00592_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\] net872 vssd1
+ vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13748__A2 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_56_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11759__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09132_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\] net858 vssd1
+ vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__and3_1
XANTENNA__09282__D1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] net907
+ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__and3_1
XANTENNA__12037__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout213_A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14173__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] vssd1 vssd1 vccd1 vccd1 net2237
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold643 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\] vssd1 vssd1 vccd1 vccd1
+ net2259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold654 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10780__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16033__A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1122_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[5\] net844 vssd1
+ vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout582_A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\] net844
+ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__and3_1
X_09896_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] net883 vssd1
+ vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__and3_1
Xhold1310 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09352__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1332 _02127_ vssd1 vssd1 vccd1 vccd1 net2948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1343 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\] net879
+ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__and3_1
Xhold1354 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2970 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout847_A _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1365 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1387 _03493_ vssd1 vssd1 vccd1 vccd1 net3003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12500__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__o21a_1
Xhold1398 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold258_A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09081__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08917__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__B _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10740_ net545 _06953_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__and2_2
XFILLER_0_138_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16976__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _06778_ _06832_ _06933_ _06934_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__or4_2
X_12410_ net2454 net225 net421 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13390_ net2563 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1
+ vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09748__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08652__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ net2360 net198 net490 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16206__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ net1239 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
X_12272_ net2668 net236 net431 vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__mux2_1
X_14011_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\] _04149_ _04191_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\] vssd1 vssd1 vccd1 vccd1 _04192_
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_120_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11223_ _05823_ net337 vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18034__1600 vssd1 vssd1 vccd1 vccd1 net1600 _18034__1600/LO sky130_fd_sc_hd__conb_1
XFILLER_0_43_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11154_ net544 _07271_ _07417_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\] net899 vssd1
+ vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15782__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15962_ net1336 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__inv_2
X_11085_ _06179_ _06601_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__and2_1
XANTENNA__13675__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17701_ clknet_leaf_72_wb_clk_i _03261_ _01540_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10036_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[4\] net873 vssd1
+ vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__and3_1
X_14913_ net1287 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ net1354 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__inv_2
XANTENNA__14398__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ clknet_leaf_142_wb_clk_i _03192_ _01495_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_18049__1611 vssd1 vssd1 vccd1 vccd1 net1611 _18049__1611/LO sky130_fd_sc_hd__conb_1
XANTENNA__11815__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12410__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14844_ net1357 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
XANTENNA__08396__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17563_ clknet_leaf_36_wb_clk_i _03123_ _01426_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11534__B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14775_ net1326 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11987_ net3007 net249 net470 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ clknet_leaf_102_wb_clk_i net1905 _00377_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13726_ _04464_ _04019_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17494_ clknet_leaf_33_wb_clk_i _03054_ _01357_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ _06910_ _07201_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ clknet_leaf_81_wb_clk_i _02073_ _00308_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13657_ _03772_ _03792_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__xor2_1
X_10869_ net526 _07059_ _07132_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12608_ net2154 net223 net396 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16376_ clknet_leaf_110_wb_clk_i net1787 _00244_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13588_ net189 _07922_ _03928_ net768 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__o211a_1
XANTENNA__09803__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12365__B _07835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18115_ net1489 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15327_ net1296 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ net3125 net287 net403 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14155__A2 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18046_ net1608 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15258_ net1265 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13363__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14209_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\] _04253_ _04276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\]
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__a221o_1
XANTENNA__13477__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15189_ net1174 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11709__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 _03562_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_4
Xfanout419 net422 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_6
XANTENNA__09393__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__B _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_103_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08790__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] net635 _05997_
+ _05999_ _06011_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__a2111o_1
XANTENNA__16849__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[23\] net735 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22o_1
X_09681_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\] net909 vssd1
+ vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13924__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[29\] net659 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\]
+ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a221o_1
XANTENNA__11725__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08563_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13969__A2 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ net1003 net885 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__and2_1
XANTENNA__10101__B1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout428_A _08024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11460__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09568__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] net576 net577 vssd1 vssd1
+ vccd1 vccd1 _05379_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12990__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1337_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09046_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] net576 net577 vssd1 vssd1
+ vccd1 vccd1 _05310_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout797_A team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold440 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] vssd1 vssd1 vccd1 vccd1
+ net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold451 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold462 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold473 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[22\] vssd1 vssd1 vccd1 vccd1
+ net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_4
Xfanout931 _04663_ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_4
XANTENNA__08781__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09948_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net591 vssd1 vssd1 vccd1
+ vccd1 _06212_ sky130_fd_sc_hd__and2_1
Xfanout942 _04655_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17774__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout953 net955 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10242__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_2
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11668__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09879_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] net667 vssd1 vssd1
+ vccd1 vccd1 _06143_ sky130_fd_sc_hd__or2_1
XANTENNA__12865__C1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 net998 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1151 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ net2222 net227 net475 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__mux2_1
XANTENNA__12230__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 team_01_WB.instance_to_wrap.cpu.f0.num\[19\] vssd1 vssd1 vccd1 vccd1 net2789
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ net3145 net607 net589 _03596_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
Xhold1184 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08647__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ net778 _07959_ _07960_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14560_ net1332 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
X_11772_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\] net674 net777 vssd1 vssd1
+ vccd1 vccd1 _07905_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13511_ _03758_ _03862_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10723_ _06860_ _06862_ _06865_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11840__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14491_ net1358 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16230_ clknet_leaf_37_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[11\]
+ _00098_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13442_ net1116 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] net781 vssd1 vssd1
+ vccd1 vccd1 _03795_ sky130_fd_sc_hd__and3_1
X_10654_ _06902_ _06917_ _06911_ _06908_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18106__1480 vssd1 vssd1 vccd1 vccd1 _18106__1480/HI net1480 sky130_fd_sc_hd__conb_1
XFILLER_0_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13373_ net3193 net328 net352 net1874 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
X_16161_ clknet_leaf_90_wb_clk_i _01829_ _00029_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15777__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10585_ _06845_ _06848_ _04716_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ net1208 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
XANTENNA__14137__A2 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ net2123 net245 net429 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
XANTENNA__09775__A _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16092_ net1403 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13345__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ net1907 net262 net437 vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__mux2_1
X_15043_ net1221 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12405__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09013__A1 _05276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11206_ _07207_ _07209_ net525 vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12186_ net2925 net246 net443 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ net338 net341 _06247_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13648__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16994_ clknet_leaf_144_wb_clk_i _02554_ _00857_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ net1393 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__inv_2
XANTENNA__11659__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ _05760_ net340 net337 _05755_ _07331_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A2 _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\] net894 vssd1
+ vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12140__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ net1396 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__inv_2
XANTENNA__09015__A _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17615_ clknet_leaf_124_wb_clk_i _03175_ _01478_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14827_ net1341 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17546_ clknet_leaf_43_wb_clk_i _03106_ _01409_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14758_ net1202 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ _04558_ _04023_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17477_ clknet_leaf_135_wb_clk_i _03037_ _01340_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14689_ net1402 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16428_ clknet_leaf_103_wb_clk_i _02056_ _00291_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16521__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16359_ clknet_leaf_76_wb_clk_i _01993_ _00227_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14128__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13336__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18029_ net1423 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_23_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17797__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16671__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout205 _07888_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout216 _07943_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout227 _07911_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlymetal6s2s_1
X_09802_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\] net722 net713 _06064_
+ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__a2111o_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
Xfanout249 _07953_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10062__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09733_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\] net878
+ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09851__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout280_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08515__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13146__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[11\] net844
+ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__and3_1
XANTENNA__10322__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] net734 net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a22o_1
X_09595_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] net845 vssd1
+ vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout545_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08546_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\] net930 vssd1
+ vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08764__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ net1075 net893 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__and2_4
XANTENNA_fanout712_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08483__B net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09298__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15597__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13575__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10389__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10237__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10928__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10370_ _06630_ _06631_ _06632_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09794__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18048__1610 vssd1 vssd1 vccd1 vccd1 net1610 _18048__1610/LO sky130_fd_sc_hd__conb_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\] net706 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12225__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ net3196 net236 net459 vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
Xhold270 _01985_ vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold281 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 _04643_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_6
XANTENNA__08939__A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_2
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_4
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_4
X_13991_ _04167_ _04178_ _04174_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a21o_1
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15730_ net1184 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
X_12942_ net1027 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1
+ vccd1 _03634_ sky130_fd_sc_hd__or2_1
XANTENNA__10313__B1 _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15661_ net1216 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
X_12873_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net1056 net366 _03583_
+ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a22o_1
X_17400_ clknet_leaf_28_wb_clk_i _02960_ _01263_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14612_ net1358 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
X_11824_ net780 _07945_ _07946_ _07947_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_16_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15592_ net1183 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12908__B _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17331_ clknet_leaf_50_wb_clk_i _02891_ _01194_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14543_ net1319 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
X_11755_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] net674 vssd1 vssd1 vccd1
+ vccd1 _07891_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17262_ clknet_leaf_55_wb_clk_i _02822_ _01125_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10706_ net534 _06953_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__and2_2
X_14474_ net1335 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
X_11686_ _07838_ _07839_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16213_ clknet_leaf_118_wb_clk_i _01880_ _00081_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_13425_ _03776_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17193_ clknet_leaf_49_wb_clk_i _02753_ _01056_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ _05622_ _06036_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__and2_1
XANTENNA__16694__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16144_ net1322 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__inv_2
XANTENNA__11041__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10568_ _06829_ _06831_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ net31 net800 net595 net1715 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__o22a_1
XANTENNA__09936__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13318__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08840__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ net2233 net286 net427 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
X_16075_ net1401 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__inv_2
XANTENNA__12135__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ net101 net814 net599 net1637 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
X_10499_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\] net657 _04759_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _06763_ sky130_fd_sc_hd__a22o_1
XANTENNA__13869__B2 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15026_ net1174 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238_ net2213 net203 net436 vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11974__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__A2 _07011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12169_ net2653 net190 net443 vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08849__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09671__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16977_ clknet_leaf_24_wb_clk_i _02537_ _00840_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_15928_ net1342 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15859_ net1188 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14586__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08400_ net1118 net929 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__and2_2
XANTENNA__13490__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09380_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\] net720 _05628_
+ _05630_ _05634_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08584__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ net3178 net2904 net1049 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ clknet_leaf_18_wb_clk_i _03089_ _01392_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08262_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\] net2787 net1039 vssd1 vssd1
+ vccd1 vccd1 _03485_ sky130_fd_sc_hd__mux2_1
XANTENNA__11280__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08193_ _04480_ _04566_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10057__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12045__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08736__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16041__A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__B1 _06805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09716_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\] net749 net737 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16567__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10520__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17812__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09647_ _05908_ _05909_ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout927_A _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08494__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] net690 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\]
+ _05827_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] net659 net608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\]
+ _04735_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a221o_1
XANTENNA__11632__B _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13260__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11124__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ net1064 _07773_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__nand2_1
XANTENNA__10074__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17962__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__A1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ net1065 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _07723_ vssd1 vssd1 vccd1
+ vccd1 _07724_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10422_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\] net735 _06672_
+ _06673_ _06674_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15120__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ net2084 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\] net818 vssd1 vssd1
+ vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
X_14190_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\] _04244_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[115\]
+ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\] net921 vssd1
+ vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and3_1
X_13141_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[93\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\]
+ net823 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13072_ net1622 net836 net356 _03701_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XANTENNA__09519__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\] net910 vssd1
+ vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__o21a_1
XANTENNA__11326__A2 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net3102 net262 net464 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_1
X_16900_ clknet_leaf_139_wb_clk_i _02460_ _00763_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08727__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17342__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ clknet_leaf_99_wb_clk_i net2359 _01700_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10534__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ clknet_leaf_1_wb_clk_i _02391_ _00694_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout580 _04722_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
Xfanout591 _04848_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_2
X_16762_ clknet_leaf_34_wb_clk_i _02322_ _00625_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13974_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[3\] net584 vssd1 vssd1
+ vccd1 vccd1 _04165_ sky130_fd_sc_hd__or2_1
XANTENNA__13484__C1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15713_ net1313 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17492__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__S1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ team_01_WB.instance_to_wrap.a1.ADR_I\[17\] net604 net586 _03621_ vssd1 vssd1
+ vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16693_ clknet_leaf_24_wb_clk_i _02253_ _00556_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15644_ net1279 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ net2182 net311 net369 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13787__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net776 _07931_ _07932_ _07933_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15575_ net1239 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09455__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12787_ net2273 net245 net377 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17314_ clknet_leaf_0_wb_clk_i _02874_ _01177_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14526_ net1323 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11738_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] net674 vssd1 vssd1 vccd1
+ vccd1 _07877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11969__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17245_ clknet_leaf_129_wb_clk_i _02805_ _01108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14457_ net1391 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XANTENNA__10873__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11669_ net1819 net1159 net569 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1
+ vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15030__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18129__1503 vssd1 vssd1 vccd1 vccd1 _18129__1503/HI net1503 sky130_fd_sc_hd__conb_1
X_13408_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _06717_ vssd1 vssd1
+ vccd1 vccd1 _03761_ sky130_fd_sc_hd__and2_1
XANTENNA__09758__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17176_ clknet_leaf_30_wb_clk_i _02736_ _01039_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08343__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388_ net1328 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16127_ net1398 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13339_ net18 net801 net596 net2582 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09963__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16058_ net1405 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08718__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15009_ net1291 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] net918
+ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11717__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17835__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] net937 vssd1
+ vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13932__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09694__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] net920
+ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17985__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09203__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09363_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\] net961 vssd1
+ vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08314_ net2747 net2695 net1047 vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11253__A1 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ net978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[14\] net943 vssd1
+ vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__and3_1
XANTENNA__11253__B2 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08245_ net2205 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10783__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout410_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1152_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08176_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] _04566_ _04577_ vssd1 vssd1 vccd1
+ vccd1 _04578_ sky130_fd_sc_hd__a21o_1
XANTENNA__09749__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08253__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10764__A0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XANTENNA__12503__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _05345_ net334 net332 _05346_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12710_ net1984 net254 net383 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10295__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13690_ team_01_WB.instance_to_wrap.a1.curr_state\[0\] _03741_ _04011_ vssd1 vssd1
+ vccd1 vccd1 _04013_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12641_ net2711 net223 net393 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10047__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15360_ net1286 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
X_12572_ net2674 net289 net399 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__mux2_1
XANTENNA__08952__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] _04450_ net1366 vssd1
+ vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11795__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ net483 _07761_ net319 vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15291_ net1317 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08660__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17708__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17030_ clknet_leaf_136_wb_clk_i _02590_ _00893_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14242_ _04153_ _04393_ _04395_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__or4_1
X_11454_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] _07706_ vssd1 vssd1 vccd1 vccd1
+ _07707_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10706__B _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] net917
+ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__and3_1
X_14173_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\] _04249_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\]
+ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__a221o_1
X_11385_ net525 _07592_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ net3008 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\] net819 vssd1 vssd1
+ vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XANTENNA__09783__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10336_ _06211_ _06245_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17858__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\] net909 vssd1
+ vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__and3_1
XANTENNA__12413__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13055_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\] _03689_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__mux2_1
X_17932_ clknet_leaf_81_wb_clk_i net1792 _01752_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08176__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1320 net1321 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ net2737 net205 net465 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
XANTENNA__09373__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1331 net1333 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17863_ clknet_leaf_102_wb_clk_i net2553 _01683_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10198_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] net937 vssd1
+ vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__and3_1
Xfanout1342 net1349 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__buf_4
Xfanout1353 net1360 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__clkbuf_4
Xfanout1364 net1365 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__buf_4
Xfanout1375 net1376 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__buf_4
XANTENNA__16882__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16814_ clknet_leaf_52_wb_clk_i _02374_ _00677_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_17794_ clknet_leaf_70_wb_clk_i _03351_ _01615_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout1386 net1387 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__buf_4
XFILLER_0_17_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1397 net1398 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__buf_2
XANTENNA__10160__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16745_ clknet_leaf_38_wb_clk_i _02305_ _00608_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13957_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\] _04149_ vssd1 vssd1
+ vccd1 vccd1 _04150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11483__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12908_ net1025 _07196_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__nand2_1
X_16676_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[30\]
+ _00539_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ net2370 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09023__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15627_ net1211 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
X_12839_ net2342 net225 net370 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09958__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15558_ net1274 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14509_ net1344 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XANTENNA__12983__B2 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17388__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ net1288 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08030_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] vssd1 vssd1 vccd1 vccd1 _04461_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_114_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17228_ clknet_leaf_44_wb_clk_i _02788_ _01091_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
Xinput41 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
XFILLER_0_126_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09396__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput52 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold803 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput74 wbs_we_i vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
Xhold814 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ clknet_leaf_121_wb_clk_i _02719_ _01022_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold825 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\] vssd1 vssd1 vccd1 vccd1
+ net2441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold847 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold858 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _06212_ _06244_ net582 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__mux2_4
Xhold869 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08801__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08932_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\] net632 net629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a22o_1
XANTENNA__12323__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08167__B2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1503 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\] vssd1 vssd1 vccd1 vccd1
+ net3119 sky130_fd_sc_hd__dlygate4sd3_1
X_08863_ _05123_ _05124_ _05125_ _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout193_A _07874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1514 _02135_ vssd1 vssd1 vccd1 vccd1 net3130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1536 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1547 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08794_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] net628 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a22o_1
Xhold1569 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10778__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout360_A _03665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A _08016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] net662 _05656_
+ _05661_ _05670_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12993__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout625_A _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14774__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09346_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] net620 _05594_
+ _05599_ _05601_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_34_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11777__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] net644 _05516_
+ _05519_ _05526_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10807__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08491__B net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14176__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08228_ net1708 net784 _00020_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16755__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout994_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08159_ net1742 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1
+ vccd1 vccd1 _03536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ _06277_ _06347_ net505 vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ _06347_ _06382_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08158__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10052_ _06277_ net547 vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__nand2_1
XANTENNA__10261__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ net1342 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09107__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ net486 net564 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1
+ vccd1 _04109_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14100__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18128__1502 vssd1 vssd1 vccd1 vccd1 _18128__1502/HI net1502 sky130_fd_sc_hd__conb_1
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09658__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ net1326 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16530_ clknet_leaf_64_wb_clk_i _02158_ _00393_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13742_ _07720_ _07773_ _04017_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a21bo_1
X_10954_ _07214_ _07216_ _07217_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08385__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16461_ clknet_leaf_80_wb_clk_i net2980 _00324_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_13673_ _07991_ _03998_ net187 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__mux2_1
X_10885_ net527 _07053_ _06971_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18200_ net1574 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
XANTENNA__17530__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15412_ net1244 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
X_12624_ net2807 net260 net398 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
X_16392_ clknet_leaf_72_wb_clk_i _02020_ _00255_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_112_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ net1505 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
XANTENNA__12916__B _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12965__B2 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15343_ net1200 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
X_12555_ net3158 net315 net404 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12408__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11506_ net1062 _07732_ _07749_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__or3_1
X_18062_ net1436 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_41_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10440__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15274_ net1196 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
X_12486_ net2070 net268 net413 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
X_17013_ clknet_leaf_8_wb_clk_i _02573_ _00876_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ _04375_ _04377_ _04379_ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__or4_1
X_11437_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] net1162 _04596_ _07683_ vssd1
+ vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10155__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13390__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14156_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\] _04260_ _04275_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\]
+ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11368_ net332 _07630_ _07631_ _04958_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13107_ net1964 net837 net357 _03723_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a22o_1
X_10319_ _06579_ _06580_ _06581_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12143__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14087_ _04226_ net787 _04236_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__and3_4
X_11299_ _06029_ _07498_ _05963_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08149__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_119_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13038_ net1694 net835 net355 _03678_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
XANTENNA__09018__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17915_ clknet_leaf_82_wb_clk_i net2020 _01735_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11982__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1
+ net1150 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1161 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 net1161
+ sky130_fd_sc_hd__buf_4
XFILLER_0_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17846_ clknet_leaf_89_wb_clk_i _03396_ _01666_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout1172 _00026_ vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_4
Xfanout1183 net1185 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__buf_4
XANTENNA__08857__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1194 net1302 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17060__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14989_ net1212 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
X_17777_ clknet_leaf_105_wb_clk_i _03335_ _01598_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16628__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10259__A2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16728_ clknet_leaf_27_wb_clk_i _02288_ _00591_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11197__A2_N _06382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659_ clknet_leaf_96_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[13\]
+ _00522_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14594__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09200_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\] net878
+ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08592__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12956__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09131_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\] net873 vssd1
+ vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__and3_1
XANTENNA__08624__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11222__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[18\] net877
+ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_96_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold600 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout206_A _07879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold611 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\] vssd1 vssd1 vccd1 vccd1 net2227
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10065__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09585__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold644 team_01_WB.instance_to_wrap.a1.ADR_I\[18\] vssd1 vssd1 vccd1 vccd1 net2260
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09854__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold655 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold677 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09964_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] net887 vssd1
+ vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__and3_1
XANTENNA__12053__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold699 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\] vssd1 vssd1 vccd1 vccd1
+ net2315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16158__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08915_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\] net898 vssd1
+ vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__and3_1
XANTENNA__17403__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[6\] net905 vssd1
+ vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__and3_1
XANTENNA__12988__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1300 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 team_01_WB.instance_to_wrap.cpu.f0.state\[0\] vssd1 vssd1 vccd1 vccd1 net2927
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10498__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] net871
+ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__and3_1
Xhold1333 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12892__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1344 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1366 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1377 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\] vssd1 vssd1 vccd1 vccd1
+ net2993 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout742_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08777_ _05033_ _05034_ _05038_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__or4_4
Xhold1388 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[73\] vssd1 vssd1 vccd1 vccd1
+ net3004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\] vssd1 vssd1 vccd1 vccd1
+ net3015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17553__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09598__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10670_ _06668_ _06721_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09329_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\] net903
+ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__and3_1
XANTENNA__12947__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12228__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14149__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10422__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ net2782 net289 net490 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ net3245 net204 net433 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[4\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__or4_1
XANTENNA__09576__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13372__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11222_ _07253_ _07256_ net541 vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09040__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _06319_ net341 _07416_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17083__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[3\] net853 vssd1
+ vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__and3_1
X_15961_ net1330 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__inv_2
X_11084_ _06178_ _06896_ _07346_ net324 vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12898__S net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14679__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17700_ clknet_leaf_72_wb_clk_i _03260_ _01539_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10035_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\] net848 vssd1
+ vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__and3_1
X_14912_ net1273 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
X_15892_ net1350 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ net1384 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
X_17631_ clknet_leaf_2_wb_clk_i _03191_ _01494_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08396__B net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17562_ clknet_leaf_34_wb_clk_i _03122_ _01425_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ net1307 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
X_11986_ net1925 net276 net470 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16513_ clknet_leaf_99_wb_clk_i _02141_ _00376_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ sky130_fd_sc_hd__dfstp_1
X_13725_ _07681_ _04041_ _04043_ net783 net1630 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o32a_1
XANTENNA__16920__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17493_ clknet_leaf_25_wb_clk_i _03053_ _01356_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10937_ _06907_ _07200_ _05622_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_58_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12927__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16444_ clknet_leaf_107_wb_clk_i net1903 _00307_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_13656_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _03985_ net1067 vssd1
+ vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__mux2_1
X_10868_ net526 _07131_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12938__A1 _07551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09301__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ net2346 net228 net395 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XANTENNA__08843__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16375_ clknet_leaf_111_wb_clk_i net1954 _00243_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08606__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12138__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ net189 _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10799_ _04883_ _04828_ net501 vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__mux2_1
X_18114_ net1488 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12365__C _07840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15326_ net1312 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ net2888 net232 net405 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11977__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18045_ net1607 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_15257_ net1192 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
X_12469_ net2744 net238 net411 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XANTENNA__16134__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14208_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\] _04238_ _04242_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\]
+ _04363_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__a221o_1
XANTENNA__13363__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17426__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net1242 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XANTENNA__09031__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] _04229_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[113\]
+ _04290_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a221o_1
Xfanout409 _03562_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09319__B1 _05581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16450__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] net950
+ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09680_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\] net905
+ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__and3_1
XANTENNA__12601__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_143_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08631_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\] net639 net615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a22o_1
X_17829_ clknet_leaf_89_wb_clk_i _03386_ _01650_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ _04815_ _04817_ _04822_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__or4_4
XFILLER_0_72_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09098__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ net1018 net858 vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__and2_2
XFILLER_0_33_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09849__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12929__A1 team_01_WB.instance_to_wrap.a1.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08753__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout323_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] net762 _05376_ _05377_
+ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09045_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] net760 _05307_ _05308_
+ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a22o_4
XFILLER_0_130_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1232_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18127__1501 vssd1 vssd1 vccd1 vccd1 _18127__1501/HI net1501 sky130_fd_sc_hd__conb_1
XFILLER_0_103_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13354__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold430 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08261__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold441 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold485 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\] vssd1 vssd1 vccd1 vccd1
+ net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13106__A1 _06381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold496 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout910 net912 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10523__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09881__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout921 net923 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
X_09947_ _06209_ _06210_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] net761
+ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a2bb2o_4
Xfanout943 _04655_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout957_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout976 net993 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09878_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net579 net591 vssd1 vssd1
+ vccd1 vccd1 _06142_ sky130_fd_sc_hd__and3_1
Xfanout987 net991 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11668__B2 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08497__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1152 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _05082_ _05090_ _05091_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__or4_1
XANTENNA__16943__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\] vssd1 vssd1 vccd1 vccd1
+ net2779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\] vssd1 vssd1 vccd1 vccd1
+ net2801 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11127__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1196 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\] vssd1 vssd1 vccd1 vccd1
+ net2812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11840_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\] net679 net780 vssd1 vssd1
+ vccd1 vccd1 _07961_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11771_ net675 _07611_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13290__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _03758_ _03759_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10722_ _04797_ net338 net336 _04796_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_95_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14490_ net1358 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09121__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] net1156 net765 vssd1 vssd1
+ vccd1 vccd1 _03794_ sky130_fd_sc_hd__and3_1
X_10653_ _06903_ _06914_ _06916_ _05963_ _06915_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__a221o_1
XANTENNA__14962__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16160_ clknet_leaf_90_wb_clk_i _01828_ _00028_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13372_ net2677 net328 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1
+ vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17449__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08960__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10584_ _04486_ net1155 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _06846_ vssd1
+ vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11797__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15111_ net1197 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
X_12323_ net2975 net314 net428 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16091_ net1400 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__inv_2
XANTENNA__13345__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15042_ net1267 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
X_12254_ net2210 net268 net438 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ net539 _07465_ _07468_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12185_ net2498 net276 net444 vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09791__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ _06245_ net335 vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13648__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16993_ clknet_leaf_135_wb_clk_i _02553_ _00856_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13517__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ net1395 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__inv_2
XANTENNA__12421__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11659__B2 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _05753_ _06985_ net331 _05759_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A3 _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[4\] net859 vssd1
+ vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__and3_1
XANTENNA__08838__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15875_ net1393 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17614_ clknet_leaf_53_wb_clk_i _03174_ _01477_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14826_ net1341 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14073__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ net1228 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
X_17545_ clknet_leaf_49_wb_clk_i _03105_ _01408_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13281__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ net2588 net195 net469 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09485__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08827__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13708_ net1061 net485 _04028_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1
+ vccd1 vccd1 _04030_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17476_ clknet_leaf_139_wb_clk_i _03036_ _01339_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14688_ net1405 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XANTENNA__08346__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09669__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16427_ clknet_leaf_100_wb_clk_i _02055_ _00290_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_13639_ _03799_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16358_ clknet_leaf_85_wb_clk_i _01992_ _00226_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09966__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15309_ net1214 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16289_ clknet_leaf_85_wb_clk_i _01923_ _00157_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16816__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18028_ net1422 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09004__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout206 _07879_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[7\] net728 _06046_ _06054_
+ _06055_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a2111o_1
Xfanout217 _07943_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
Xfanout228 _07911_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
Xfanout239 net241 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\] _04750_
+ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__and3_1
XANTENNA__11736__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11455__B team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09663_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\] net911
+ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout273_A _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\] net750 net719 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a22o_1
X_09594_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\] net871 vssd1
+ vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08545_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\] net956 vssd1
+ vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout440_A _08021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13162__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ net1003 net903 vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__and2_4
XFILLER_0_18_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout705_A _04681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10518__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13575__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09243__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11050__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16496__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12506__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09028_ net978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] net940 vssd1
+ vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold260 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[30\] vssd1 vssd1 vccd1 vccd1
+ net1876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17891__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_6
Xfanout751 _04641_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12241__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout762 _04636_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_4
X_13990_ _04175_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__xor2_1
Xfanout773 _04625_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
Xfanout784 _04512_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_4
Xfanout795 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1 vccd1 net795
+ sky130_fd_sc_hd__buf_2
X_12941_ net1026 _07344_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15660_ net1251 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12872_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] _07023_ net1025 vssd1 vssd1
+ vccd1 vccd1 _03583_ sky130_fd_sc_hd__mux2_1
XANTENNA__08955__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14611_ net1371 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11823_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\] net676 net775 vssd1 vssd1
+ vccd1 vccd1 _07947_ sky130_fd_sc_hd__o21a_1
XANTENNA__13263__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15591_ net1195 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
X_17330_ clknet_leaf_39_wb_clk_i _02890_ _01193_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10077__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ net1323 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
X_11754_ _07863_ _07889_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09482__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17271__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ net509 _06965_ _06967_ _06968_ net527 vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__a2111o_1
X_17261_ clknet_leaf_16_wb_clk_i _02821_ _01124_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14473_ net1335 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11685_ net2369 net1169 team_01_WB.instance_to_wrap.cpu.K0.count\[0\] vssd1 vssd1
+ vccd1 vccd1 _07839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08690__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16212_ clknet_leaf_118_wb_clk_i _01879_ _00080_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _06212_ vssd1 vssd1 vccd1
+ vccd1 _03777_ sky130_fd_sc_hd__or2_1
XANTENNA__09786__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17192_ clknet_leaf_61_wb_clk_i _02752_ _01055_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ _06041_ _06043_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16143_ net1320 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08442__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ net32 net802 net596 net3091 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10567_ _06807_ _06828_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__nor2_1
XANTENNA__12416__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ net2446 net230 net429 vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ net1405 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__inv_2
X_13286_ net2059 net814 net599 net1851 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a22o_1
XANTENNA__16989__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10498_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\] net654 _04753_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[25\] _06753_ vssd1 vssd1 vccd1
+ vccd1 _06762_ sky130_fd_sc_hd__a221o_1
XANTENNA__13869__A2 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15025_ net1199 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12237_ net3056 net238 net435 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10163__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12168_ net1983 net197 net445 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XANTENNA__09952__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16219__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11119_ net339 net342 _06176_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__mux2_1
XANTENNA__12151__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ net2910 net210 net458 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
X_16976_ clknet_leaf_25_wb_clk_i _02536_ _00839_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09026__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ net1351 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__inv_2
XANTENNA__11990__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ net1188 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__inv_2
X_18126__1500 vssd1 vssd1 vccd1 vccd1 _18126__1500/HI net1500 sky130_fd_sc_hd__conb_1
XFILLER_0_133_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17614__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809_ net1384 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ net1212 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__inv_2
XANTENNA__08584__B net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08330_ net2686 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17528_ clknet_leaf_27_wb_clk_i _03088_ _01391_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09399__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08261_ net2829 net2761 net1045 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17459_ clknet_leaf_50_wb_clk_i _03019_ _01322_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08681__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09696__A _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08192_ _04579_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12326__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10791__A1 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11335__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16679__D net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11466__A team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12061__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09146__D1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09715_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\] net751 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a22o_1
XANTENNA__12996__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14777__A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout655_A _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1397_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\] net723 _04685_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09577_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] net724 _05830_ _05831_
+ _05833_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08528_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] net637 net629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\]
+ _04778_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08672__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ net781 _04715_ net681 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or3_2
XFILLER_0_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13548__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15401__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] team_01_WB.instance_to_wrap.cpu.f0.i\[4\]
+ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10421_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\] net729 net711 _06676_
+ _06679_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12236__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11140__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13140_ net2607 net2524 net819 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
X_10352_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] net931 vssd1
+ vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__and3_1
X_13071_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\] _03700_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__mux2_1
X_10283_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\] _04767_ _06544_ _06545_
+ _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13720__A1 _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ net2964 net266 net465 vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input49_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16830_ clknet_leaf_3_wb_clk_i _02390_ _00693_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_2
XANTENNA__14276__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_4
Xfanout592 _04848_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_1
X_13973_ _03554_ _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__or2_1
X_16761_ clknet_leaf_125_wb_clk_i _02321_ _00624_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14687__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12924_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] net1053 net364 _03620_
+ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__a22o_1
X_15712_ net1289 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
X_16692_ clknet_leaf_12_wb_clk_i _02252_ _00555_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12039__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13236__A0 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15643_ net1298 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
X_12855_ net1841 net259 net369 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17787__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ net681 _07265_ net776 vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15574_ net1305 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12786_ net2871 net314 net375 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14525_ net1322 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17313_ clknet_leaf_136_wb_clk_i _02873_ _01176_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11737_ _07865_ _07875_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08663__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10158__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14456_ net1390 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17244_ clknet_leaf_13_wb_clk_i _02804_ _01107_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17017__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09207__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ net3023 net1160 net568 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1
+ vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14200__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13407_ _03759_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08851__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ _06525_ _06880_ _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__o21ai_1
X_17175_ clknet_leaf_10_wb_clk_i _02735_ _01038_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire960 _04640_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12146__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ net1385 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
X_11599_ net496 _07814_ net2415 net838 vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_25_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16126_ net1397 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338_ net19 net799 net594 net2558 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11985__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ net1368 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__inv_2
X_13269_ net1682 net813 net599 team_01_WB.instance_to_wrap.a1.ADR_I\[22\] vssd1 vssd1
+ vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15008_ net1273 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09682__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08194__A2 _04593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__A _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14267__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16959_ clknet_leaf_2_wb_clk_i _02519_ _00822_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_09500_ net980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\] net953 vssd1
+ vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__and3_1
XANTENNA__13932__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09694__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] net956
+ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13227__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\] net935 vssd1
+ vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09446__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11789__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08313_ net3079 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09293_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] net957
+ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__and3_1
XANTENNA__08654__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout236_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08244_ net1680 net2399 net1041 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09857__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08761__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12056__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _04573_ _04574_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout403_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1145_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10764__A1 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1312_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_101_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09906__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XANTENNA__09592__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08489__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ net539 _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__nor2_1
XANTENNA__09685__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09629_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] net932 vssd1
+ vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__and3_1
XANTENNA__08893__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12640_ net3075 net229 net391 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XANTENNA__13769__B2 _00020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12571_ net2381 net233 net401 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14310_ _04450_ _04451_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15131__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ _07711_ _07739_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ net1259 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14241_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\] _04233_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\]
+ _04396_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__a221o_1
X_11453_ team_01_WB.instance_to_wrap.cpu.f0.i\[12\] net1064 _07705_ vssd1 vssd1 vccd1
+ vccd1 _07706_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _06666_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__nor2_2
X_14172_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[11\] _04252_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\]
+ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a22o_1
X_11384_ net531 _07260_ _07076_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__a21oi_1
X_13123_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\] net3129 net824 vssd1 vssd1
+ vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10335_ _06247_ _06316_ _06246_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10850__S1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13054_ _05199_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__o21a_1
X_17931_ clknet_leaf_83_wb_clk_i _03481_ _01751_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] net663 _06527_ _06528_
+ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ net2407 net238 net463 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
Xfanout1310 net1415 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_4
Xfanout1321 net1325 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1332 net1333 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__buf_4
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17862_ clknet_leaf_96_wb_clk_i _03412_ _01682_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ sky130_fd_sc_hd__dfstp_1
X_10197_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[1\] net951 vssd1
+ vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__and3_1
Xfanout1343 net1345 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__buf_4
XANTENNA__14249__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1354 net1356 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__buf_4
X_16813_ clknet_leaf_19_wb_clk_i _02373_ _00676_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1365 net1370 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__buf_2
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1376 net1379 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__buf_4
X_17793_ clknet_leaf_70_wb_clk_i _03350_ _01614_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout1387 net1388 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__buf_4
Xfanout1398 net1414 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16744_ clknet_leaf_63_wb_clk_i _02304_ _00607_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13956_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and2_1
XANTENNA__08846__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ team_01_WB.instance_to_wrap.a1.ADR_I\[22\] net606 net588 _03608_ vssd1 vssd1
+ vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
XANTENNA__11483__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16675_ clknet_leaf_112_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[29\]
+ _00538_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13887_ net2932 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_124_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12838_ net2496 net228 net367 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__mux2_1
X_15626_ net1198 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15557_ net1233 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
XANTENNA__16407__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08636__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ net2632 net231 net377 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10443__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12983__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14508_ net1361 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XANTENNA__08354__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15488_ net1286 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
XANTENNA__09677__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17227_ clknet_leaf_51_wb_clk_i _02787_ _01090_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_14439_ net1387 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_1
XFILLER_0_128_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput42 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput64 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16557__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold804 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ clknet_leaf_140_wb_clk_i _02718_ _01021_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold815 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[27\] vssd1 vssd1 vccd1 vccd1
+ net2431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold826 _02106_ vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17802__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold837 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ net1363 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__inv_2
X_09980_ _06240_ _06242_ _06243_ _06213_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__o31a_4
X_17089_ clknet_leaf_137_wb_clk_i _02649_ _00952_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12604__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold859 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08931_ _05191_ _05192_ _05193_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10632__B _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08862_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\] net656 _05110_
+ _05112_ _05120_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1504 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\] vssd1 vssd1 vccd1 vccd1
+ net3120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1526 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1537 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3153 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13448__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08793_ _05053_ _05054_ _05055_ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1548 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\] vssd1 vssd1 vccd1 vccd1
+ net3175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09116__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15216__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08875__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\] net644 _05658_
+ _05660_ _05662_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09419__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09345_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\] net616 _05589_ _05598_
+ _05604_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08627__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13170__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10434__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09276_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\] net633 _05527_
+ _05536_ _05538_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08227_ net785 net486 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__or2_2
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10095__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09884__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ net1737 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1
+ vccd1 vccd1 _03537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17482__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout987_A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08089_ _04465_ team_01_WB.instance_to_wrap.cpu.f0.num\[24\] team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ _04469_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__a22o_1
XANTENNA__12514__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10120_ _06347_ net541 vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10051_ net579 _06313_ _06279_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10969__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13810_ net2305 net784 _07681_ _04108_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ net1333 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13741_ net564 _07680_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.next_write_i
+ sky130_fd_sc_hd__or2_1
X_10953_ net321 _07021_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13672_ _03787_ _03789_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__xnor2_1
X_16460_ clknet_leaf_108_wb_clk_i _02088_ _00323_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ net520 _07046_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12623_ net2421 net299 net398 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
X_15411_ net1188 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16391_ clknet_leaf_75_wb_clk_i _02019_ _00254_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18130_ net1504 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
X_15342_ net1228 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XANTENNA__12965__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ net2760 net302 net403 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10976__A1 _07139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11505_ net483 _07749_ net319 vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__a21o_1
XANTENNA__17825__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15273_ net1205 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
X_18061_ team_01_WB.instance_to_wrap.cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net157
+ sky130_fd_sc_hd__clkbuf_1
X_12485_ net2650 net270 net411 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17012_ clknet_leaf_6_wb_clk_i _02572_ _00875_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14224_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\] _04244_ _04246_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\]
+ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a221o_1
X_11436_ _07693_ net3260 _07685_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\] _04278_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\]
+ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12424__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ net340 net338 _04957_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10733__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10823__S1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17975__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[3\] _06381_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__mux2_1
X_10318_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\] net705 _06567_ _06571_
+ _06574_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14086_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\] _04246_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[80\]
+ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a22o_1
X_11298_ net544 _07561_ _07559_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__o21a_1
X_13037_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\] _03677_ net1028 vssd1
+ vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__mux2_1
X_17914_ clknet_leaf_78_wb_clk_i _03464_ _01734_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\] net656 _06489_ _06490_
+ _06504_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10171__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1140 net1146 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1162 team_01_WB.instance_to_wrap.cpu.f0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1162 sky130_fd_sc_hd__buf_2
X_17845_ clknet_leaf_104_wb_clk_i _03395_ _01665_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09960__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1173 net1176 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_4
XANTENNA__11564__A _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1195 net1203 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
XFILLER_0_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ clknet_leaf_95_wb_clk_i _03334_ _01597_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08349__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09649__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14988_ net1263 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16727_ clknet_leaf_9_wb_clk_i _02287_ _00590_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ net1164 net1058 net3264 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[20\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__17355__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16658_ clknet_leaf_95_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[12\]
+ _00521_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08873__A _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15609_ net1191 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16589_ clknet_leaf_86_wb_clk_i _02217_ _00452_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09130_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] net887 vssd1
+ vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__and3_1
XANTENNA__12956__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__B _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] net867
+ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09200__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold601 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12334__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold645 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[114\] vssd1 vssd1 vccd1 vccd1
+ net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09963_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] net884 vssd1
+ vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] vssd1 vssd1 vccd1 vccd1
+ net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08914_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\] net905
+ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__and3_1
X_09894_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\] net908 vssd1
+ vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1010_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1108_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1312 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[20\] net863
+ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__and3_1
XANTENNA__12892__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1323 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\] vssd1 vssd1 vccd1 vccd1
+ net2939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1334 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08560__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout568_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1356 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2983 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] net721 net711 _05029_
+ _05039_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08259__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1378 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2994
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1389 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net3005 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16722__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12509__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09328_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] net861
+ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09259_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\] net910
+ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ net2613 net240 net433 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11221_ _06042_ _07483_ _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12244__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14025__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _06316_ _06983_ net331 _06317_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__o22a_1
XANTENNA__09119__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] net894 vssd1
+ vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13864__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15960_ net1330 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__inv_2
X_11083_ _06896_ _07346_ _06178_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08958__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ net1294 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
X_10034_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\] net908 vssd1
+ vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__and3_1
X_15891_ net1350 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__inv_2
XANTENNA__16252__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ clknet_leaf_3_wb_clk_i _03190_ _01493_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ net1384 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
X_18085__1459 vssd1 vssd1 vccd1 vccd1 _18085__1459/HI net1459 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17561_ clknet_leaf_18_wb_clk_i _03121_ _01424_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14773_ net1190 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
X_11985_ net2262 net215 net470 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16512_ clknet_leaf_103_wb_clk_i _02140_ _00375_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ sky130_fd_sc_hd__dfstp_1
X_13724_ _04027_ _04042_ net485 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09789__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ _05758_ _05760_ _07199_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__nand3_1
XANTENNA__08693__A _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17492_ clknet_leaf_4_wb_clk_i _03052_ _01355_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10110__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16443_ clknet_leaf_101_wb_clk_i net2891 _00306_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_13655_ _07379_ _03984_ net769 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__mux2_1
X_10867_ _07092_ _07095_ net509 vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__mux2_1
XANTENNA__12419__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12606_ net2655 net200 net395 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XANTENNA__13060__A1 _05276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16374_ clknet_leaf_113_wb_clk_i net1621 _00242_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
X_13586_ _03833_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ net515 _07055_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09803__A2 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18113_ net1487 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
X_15325_ net1284 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
X_12537_ net2765 net234 net403 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09020__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10166__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18044_ net1606 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15256_ net1256 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
X_12468_ net3217 net208 net413 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09955__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11559__A _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ _04503_ _04567_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__nor2_1
X_14207_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\] _04246_ _04272_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\]
+ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__a22o_1
XANTENNA__13363__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15187_ net1189 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
XANTENNA__12154__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ _07845_ _07846_ net489 vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__and3_1
XANTENNA__10177__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14138_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\] _04249_ _04261_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\]
+ _04289_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__a221o_1
XANTENNA__09319__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11993__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__and2b_1
XANTENNA__09724__D1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12874__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\] net652 net634 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\]
+ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a221o_1
X_17828_ clknet_leaf_89_wb_clk_i _03385_ _01649_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10885__B1 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[30\] net700 _04823_ _04824_
+ net711 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a2111o_1
X_17759_ clknet_leaf_80_wb_clk_i _03317_ _01580_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09699__A _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ net1107 net1111 net1114 net1108 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__and4bb_4
XANTENNA__10101__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_112_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12329__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12929__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13051__A1 _05063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[17\] net710 net758 vssd1
+ vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11469__A team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12064__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 net158 vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold442 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\] vssd1 vssd1 vccd1 vccd1
+ net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold453 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\] vssd1 vssd1 vccd1 vccd1
+ net2069 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12999__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold475 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold486 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 net2113
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13684__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08781__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] net709 net757 vssd1
+ vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17520__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net947 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_4
Xfanout955 _04642_ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_6
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_2
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_2
X_09877_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] net760 _06139_ _06140_
+ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__a22o_4
Xhold1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout852_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__B _06995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08497__B net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout988 net990 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_2
Xhold1131 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[42\] vssd1 vssd1 vccd1 vccd1
+ net2747 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout999 net1009 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] net723 _05074_ _05075_
+ _05080_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_99_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 team_01_WB.instance_to_wrap.cpu.f0.num\[18\] vssd1 vssd1 vccd1 vccd1 net2791
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 _03488_ vssd1 vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1197 _02078_ vssd1 vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\] net948
+ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__and3_1
XANTENNA__12617__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ _07861_ _07902_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10721_ _06868_ _06981_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__or2_4
XANTENNA__09402__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12239__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11840__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _03771_ _03792_ _03770_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10652_ _06027_ _05993_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13042__A1 _06772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13371_ net2037 net328 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1
+ vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ net1155 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 _06847_ sky130_fd_sc_hd__or2_4
XFILLER_0_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15110_ net1274 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
X_12322_ net2581 net304 net430 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16090_ net1394 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__inv_2
XANTENNA__17050__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15041_ net1312 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XANTENNA__13345__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net2970 net271 net435 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
XANTENNA__16618__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ net523 _07358_ _07466_ _07467_ net535 vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12184_ net2039 net215 net443 vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11135_ _07175_ _07398_ net545 vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08772__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12702__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16992_ clknet_leaf_2_wb_clk_i _02552_ _00855_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16768__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15943_ net1341 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ _07270_ _07278_ net534 vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\] net865 vssd1
+ vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ net1396 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17613_ clknet_leaf_20_wb_clk_i _03173_ _01476_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14825_ net1346 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ clknet_leaf_45_wb_clk_i _03104_ _01407_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15314__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14756_ net1183 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XANTENNA__13281__B2 team_01_WB.instance_to_wrap.a1.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11968_ net494 _08011_ _08012_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08854__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ net1061 _04028_ net485 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11292__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ _07181_ _07182_ net530 vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__mux2_1
X_17475_ clknet_leaf_133_wb_clk_i _03035_ _01338_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12149__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14687_ net1364 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11899_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16426_ clknet_leaf_107_wb_clk_i _02054_ _00289_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13033__A1 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09237__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13638_ _03802_ _03970_ _03800_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13941__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14230__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11988__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16357_ clknet_leaf_73_wb_clk_i net1643 _00225_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13569_ net767 _03911_ net966 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10398__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15308_ net1266 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16288_ clknet_leaf_86_wb_clk_i _01922_ _00156_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16298__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13336__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18027_ net1421 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XANTENNA__10193__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15239_ net1183 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout207 _07879_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlymetal6s2s_1
X_09800_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] net743 net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__a22o_1
Xfanout218 _07943_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_1
XANTENNA__10921__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 _07911_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_1
XANTENNA__12612__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13935__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09731_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\] net857 vssd1
+ vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08515__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[11\] net887 vssd1
+ vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10322__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08613_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[29\] net706 _04874_
+ _04875_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09593_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] net850 vssd1
+ vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08544_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] net944
+ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09476__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__B team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08475_ net1003 net891 vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__and2_2
XANTENNA__12059__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_A _08023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17073__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14221__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13679__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13575__A2 _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout600_A _03742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1342_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09595__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18084__1458 vssd1 vssd1 vccd1 vccd1 _18084__1458/HI net1458 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\] net962
+ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09892__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold250 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[7\] vssd1 vssd1 vccd1 vccd1
+ net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 net1877
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_01_WB.instance_to_wrap.a1.ADR_I\[12\] vssd1 vssd1 vccd1 vccd1 net1899
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold294 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12522__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 _04662_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_8
Xfanout741 _04653_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] _04666_ vssd1
+ vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__and3_1
Xfanout752 _04641_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11646__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_2
Xfanout774 net777 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_2
XFILLER_0_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10849__A0 _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_2
X_12940_ net1913 net604 net586 _03632_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
XANTENNA__10313__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12871_ _04510_ _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__nor2_2
X_14610_ net1410 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XANTENNA__15134__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ net679 _07535_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__nand2_1
X_15590_ net1287 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17416__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09132__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14541_ net1319 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11753_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _07862_ vssd1 vssd1
+ vccd1 vccd1 _07889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10704_ net509 net501 _04828_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_51_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17260_ clknet_leaf_44_wb_clk_i _02820_ _01123_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ net2844 _07838_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__xor2_1
X_14472_ net1336 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08690__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14212__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16211_ clknet_leaf_117_wb_clk_i _01878_ _00079_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ _06319_ _06887_ _06890_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__a31o_2
X_13423_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ net592 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17191_ clknet_leaf_131_wb_clk_i _02751_ _01054_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16440__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17566__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16142_ net1320 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13354_ net33 net799 net594 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1
+ vccd1 vccd1 _01926_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10566_ _06807_ _06828_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12305_ net2536 net234 net427 vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
XANTENNA__13318__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13285_ net103 net813 net599 net1623 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
X_16073_ net1376 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__inv_2
X_10497_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] net659 net608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\]
+ _06760_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12236_ net3065 net207 net436 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
X_15024_ net1250 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16590__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08745__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11837__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15309__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ net494 _08008_ _08017_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14279__B1 net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ _06175_ net335 vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__and2_1
XANTENNA__08849__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12098_ net3228 net292 net456 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__mux2_1
X_16975_ clknet_leaf_54_wb_clk_i _02535_ _00838_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11049_ _06828_ net334 net332 _06831_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__o2bb2a_1
X_15926_ net1351 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11501__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XANTENNA__09170__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ net1246 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11572__A team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14808_ net1384 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15788_ net1265 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__inv_2
X_17527_ clknet_leaf_11_wb_clk_i _03087_ _01390_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14739_ net1323 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08130__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17909__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ net2735 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\] net1045 vssd1 vssd1
+ vccd1 vccd1 _03487_ sky130_fd_sc_hd__mux2_1
X_17458_ clknet_leaf_39_wb_clk_i _03018_ _01321_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13006__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08881__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14203__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16409_ clknet_leaf_86_wb_clk_i _02037_ _00272_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ sky130_fd_sc_hd__dfstp_1
X_08191_ _04586_ _04588_ _04590_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__or4_2
XFILLER_0_85_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17389_ clknet_leaf_21_wb_clk_i _02949_ _01252_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12607__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16933__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10354__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08736__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12342__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14123__A _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\] net953 vssd1
+ vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17439__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09645_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\] net728 _05896_
+ _05902_ _05904_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1292_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11482__A _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09576_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[8\] net721 net711 _05826_
+ _05832_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09449__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08527_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] net655 net617 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[31\]
+ _04779_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a221o_1
XANTENNA__13796__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout815_A _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09887__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ net764 _04719_ _04720_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12517__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ net985 net945 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10420_ _06677_ _06681_ _06682_ _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ _06607_ _06612_ _05212_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10264__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13070_ _05480_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__o21a_1
X_10282_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] net906 vssd1
+ vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12021_ net2167 net271 net463 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08727__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10534__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09127__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14968__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 _07804_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_2
X_16760_ clknet_leaf_28_wb_clk_i _02320_ _00623_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_4
X_13972_ _04163_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__inv_2
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11796__A1_N net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15711_ net1294 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
X_12923_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] _07265_ net1027 vssd1 vssd1
+ vccd1 vccd1 _03620_ sky130_fd_sc_hd__mux2_1
X_16691_ clknet_leaf_55_wb_clk_i _02251_ _00554_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11392__A _07243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16806__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15642_ net1267 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
X_12854_ net2171 net298 net369 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18199__1573 vssd1 vssd1 vccd1 vccd1 _18199__1573/HI net1573 sky130_fd_sc_hd__conb_1
X_11805_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] net676 vssd1 vssd1 vccd1
+ vccd1 _07932_ sky130_fd_sc_hd__or2_1
XANTENNA__11247__B1 _06870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15573_ net1173 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12785_ net1986 net304 net375 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17312_ clknet_leaf_2_wb_clk_i _02872_ _01175_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14524_ net1409 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
X_11736_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _07864_ vssd1 vssd1
+ vccd1 vccd1 _07875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17243_ clknet_leaf_37_wb_clk_i _02803_ _01106_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14455_ net1390 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12427__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ net1745 net1160 net568 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1
+ vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _06663_ vssd1 vssd1
+ vccd1 vccd1 _03759_ sky130_fd_sc_hd__nand2_1
X_17174_ clknet_leaf_30_wb_clk_i _02734_ _01037_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10618_ _06485_ net517 vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11598_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[27\] net572 vssd1 vssd1 vccd1
+ vccd1 _07814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14386_ net1352 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08966__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16125_ net1394 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10549_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\] net660 net631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\]
+ _06812_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a221o_1
X_13337_ net20 net801 net596 net2923 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10174__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ net1374 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__inv_2
XANTENNA__09963__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ net90 net816 net600 net1618 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a22o_1
X_15007_ net1298 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08718__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12162__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ net2580 net248 net439 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13199_ net2149 net2128 net830 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10190__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16958_ clknet_leaf_12_wb_clk_i _02518_ _00821_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08876__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09143__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ net1341 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__inv_2
XANTENNA__08351__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16889_ clknet_leaf_125_wb_clk_i _02449_ _00752_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_18083__1457 vssd1 vssd1 vccd1 vccd1 _18083__1457/HI net1457 sky130_fd_sc_hd__conb_1
X_09430_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] net953
+ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09361_ net1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[13\] net913
+ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__and3_1
XANTENNA__09203__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08312_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[44\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09292_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\] net949 vssd1
+ vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_12 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ net2861 net2859 net1048 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__mux2_1
XANTENNA__09500__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17881__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12337__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _07911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _04570_ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17111__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11961__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1138_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_101_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XANTENNA__12072__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1305_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16829__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ _05823_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09559_ _05788_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12570_ net3147 net235 net399 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08952__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10452__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07745_ _07758_ _07760_ vssd1
+ vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12247__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11452_ _04475_ _07704_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nor2_2
XFILLER_0_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14240_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] _04256_ _04278_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[38\]
+ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10403_ _06643_ _06664_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__nor2_1
X_14171_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] _04264_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[11\]
+ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a221o_1
X_11383_ _07004_ _07486_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__nand2_1
XANTENNA_input61_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _06319_ _06597_ _06316_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__o21a_1
X_13122_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[112\] net1889 net819 vssd1 vssd1
+ vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09783__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17604__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17930_ clknet_leaf_78_wb_clk_i _03480_ _01750_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_13053_ net3202 net835 net356 _03688_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10265_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\] net869 vssd1
+ vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1300 net1301 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__clkbuf_4
X_12004_ net2828 net208 net465 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__mux2_1
Xfanout1311 net1313 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17861_ clknet_leaf_104_wb_clk_i _03411_ _01681_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09373__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1322 net1324 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__buf_4
X_10196_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] net922 vssd1
+ vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1333 net1337 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__clkbuf_4
Xfanout1344 net1345 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__buf_4
X_16812_ clknet_leaf_45_wb_clk_i _02372_ _00675_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1355 net1356 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__buf_4
Xfanout1366 net1370 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12710__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17792_ clknet_leaf_70_wb_clk_i _03349_ _01613_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08696__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1377 net1379 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__buf_4
Xfanout390 _03567_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_4
Xfanout1388 net1389 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__clkbuf_4
Xfanout1399 net1400 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__buf_4
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16743_ clknet_leaf_126_wb_clk_i _02303_ _00606_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13955_ _04509_ _04146_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12906_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] net1055 net365 _03607_
+ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16674_ clknet_leaf_114_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[28\]
+ _00537_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10140__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ team_01_WB.EN_VAL_REG net601 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__or2_1
XFILLER_0_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15625_ net1215 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ net2538 net201 net367 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
XANTENNA__09023__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10169__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12968__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ net1224 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
X_12768_ net2981 net236 net375 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09958__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14507_ net1344 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XANTENNA__12157__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ _07859_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15487_ net1295 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10466__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12699_ net2968 net206 net385 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17226_ clknet_leaf_41_wb_clk_i _02786_ _01089_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14438_ net1395 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
Xinput43 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11996__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput54 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
X_17157_ clknet_leaf_135_wb_clk_i _02717_ _01020_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput65 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14369_ net1326 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
Xhold805 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold816 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ net1403 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_137_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17284__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold838 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ clknet_leaf_142_wb_clk_i _02648_ _00951_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold849 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16039_ net1368 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__inv_2
X_08930_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] net657 _05173_
+ _05175_ _05177_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09990__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\] net614 _05102_
+ _05113_ _05117_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08572__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1505 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[55\] vssd1 vssd1 vccd1 vccd1
+ net3121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 team_01_WB.instance_to_wrap.cpu.K0.code\[0\] vssd1 vssd1 vccd1 vccd1 net3143
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12620__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13448__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08792_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\] net637 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a22o_1
Xhold1538 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1549 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\] vssd1 vssd1 vccd1 vccd1
+ net3165 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11744__B _07640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10682__A1 _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\] net612 _05665_ _05666_
+ _05667_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout346_A _06869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1088_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09344_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\] net609 _05588_
+ _05600_ _05605_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_34_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09230__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\] net631 _05524_
+ _05525_ _05533_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout513_A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_136_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08226_ _04502_ net1161 team_01_WB.instance_to_wrap.cpu.f0.state\[7\] _04620_ vssd1
+ vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14176__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16501__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17627__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ net1689 net552 net349 net1063 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08088_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] team_01_WB.instance_to_wrap.cpu.f0.num\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout882_A _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18198__1572 vssd1 vssd1 vccd1 vccd1 _18198__1572/HI net1572 sky130_fd_sc_hd__conb_1
XANTENNA__17777__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ net579 _06313_ _06279_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08563__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13626__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17007__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09107__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09405__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14100__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13740_ net1763 net783 _07681_ _04055_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__o22a_1
XANTENNA__10122__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10952_ _06036_ net340 net337 _05553_ _07215_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13671_ _04501_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _03996_ _03997_
+ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10883_ _06722_ net340 net338 _06720_ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__o221a_1
X_15410_ net1175 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
X_12622_ net2038 net242 net397 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
X_16390_ clknet_leaf_75_wb_clk_i _02018_ _00253_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15341_ net1213 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12553_ net2040 net264 net404 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18060_ team_01_WB.instance_to_wrap.cpu.LCD0.lcd_en vssd1 vssd1 vccd1 vccd1 net156
+ sky130_fd_sc_hd__clkbuf_1
X_11504_ _07720_ _07739_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__nand2_1
XANTENNA__16181__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15272_ net1183 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ net2398 net248 net411 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17011_ clknet_leaf_49_wb_clk_i _02571_ _00874_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14223_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\] _04261_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\]
+ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _04592_ _07683_ _07692_ net1162 vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12705__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18082__1456 vssd1 vssd1 vccd1 vccd1 _18082__1456/HI net1456 sky130_fd_sc_hd__conb_1
X_14154_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] _04239_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__a22o_1
X_11366_ _04956_ net334 vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10733__B _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13105_ net1723 net837 net357 _03722_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
X_10317_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] net732 net714 vssd1
+ vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__a21o_1
X_14085_ net789 _04237_ _04243_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__and3_4
X_11297_ net537 _06991_ _07472_ _07560_ _07335_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__o311a_1
XFILLER_0_21_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09346__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] net654 _06492_ _06499_
+ _06506_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__a2111o_1
X_13036_ _06662_ net571 net359 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__o21a_1
X_17913_ clknet_leaf_107_wb_clk_i net2402 _01733_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09018__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1130 net1133 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_2
XANTENNA__11153__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08554__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1141 net1142 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_2
X_17844_ clknet_leaf_78_wb_clk_i _03394_ _01664_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10179_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\] net628 _06419_ _06433_
+ _06435_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12440__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1152 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1
+ net1152 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1163 net1164 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_2
Xfanout1174 net1176 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_4
Xfanout1185 net1302 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
XANTENNA__08857__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17775_ clknet_leaf_116_wb_clk_i _03333_ _01596_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1196 net1203 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_2
X_14987_ net1208 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
XANTENNA__11056__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16726_ clknet_leaf_33_wb_clk_i _02286_ _00589_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13938_ net1164 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[19\] sky130_fd_sc_hd__and3b_1
XFILLER_0_57_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657_ clknet_leaf_96_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[11\]
+ _00520_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13869_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] team_01_WB.instance_to_wrap.cpu.DM0.dhit
+ team_01_WB.instance_to_wrap.cpu.f0.state\[0\] team_01_WB.EN_VAL_REG vssd1 vssd1
+ vccd1 vccd1 _04141_ sky130_fd_sc_hd__a22o_1
XANTENNA__16148__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15608_ net1254 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16588_ clknet_leaf_72_wb_clk_i _02216_ _00451_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13602__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16524__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08592__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ net1187 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
XANTENNA__10196__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\] net881
+ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__and3_1
XANTENNA__09985__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14158__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17209_ clknet_leaf_17_wb_clk_i _02769_ _01072_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12615__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18189_ net1563 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13938__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold602 team_01_WB.instance_to_wrap.cpu.f0.num\[13\] vssd1 vssd1 vccd1 vccd1 net2218
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09585__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\] vssd1 vssd1 vccd1 vccd1
+ net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold657 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold668 _03505_ vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold679 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] net905 vssd1
+ vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08913_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\] net858 vssd1
+ vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09893_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] net873 vssd1
+ vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1302 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\] vssd1 vssd1 vccd1 vccd1
+ net2918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1313 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12350__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] net858 vssd1
+ vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12892__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1324 _03462_ vssd1 vssd1 vccd1 vccd1 net2940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 net2962
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09225__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1357 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2984 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] net727 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout463_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1379 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09879__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1372_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__A team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09598__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\] net867
+ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14149__A2 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09895__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\] net847 vssd1
+ vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13357__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08209_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] _04567_ vssd1 vssd1 vccd1 vccd1
+ _04605_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09189_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\] net896 vssd1
+ vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__and3_1
XANTENNA__12525__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _06899_ _06900_ _06912_ _06043_ net324 vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__a221o_1
XANTENNA__09576__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14025__B _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11151_ net335 _07275_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10272__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] net883 vssd1
+ vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _06892_ _07345_ _06179_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__a21o_1
XANTENNA__12868__C1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] net899 vssd1
+ vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and3_1
X_14910_ net1291 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
XANTENNA__12260__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ net1357 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09135__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ net1384 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ clknet_leaf_27_wb_clk_i _03120_ _01423_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14772_ net1256 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11984_ net2694 net278 net467 vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16511_ clknet_leaf_77_wb_clk_i _02139_ _00374_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_13723_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _04026_ vssd1 vssd1 vccd1 vccd1
+ _04042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17491_ clknet_leaf_49_wb_clk_i _03051_ _01354_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11843__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ _06899_ _06900_ _06903_ _06917_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16442_ clknet_leaf_107_wb_clk_i net2700 _00305_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13654_ _07973_ _03983_ net187 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ _06722_ _07128_ _07129_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ net2894 net286 net395 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16373_ clknet_leaf_110_wb_clk_i net1843 _00241_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09301__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _05310_ _03925_ vssd1
+ vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _06997_ _07060_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112_ net1486 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
X_15324_ net1232 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XANTENNA__15600__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\] net204 net405 vssd1
+ vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13348__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18043_ net1605 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15255_ net1243 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
X_12467_ net2799 net190 net411 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XANTENNA__12435__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\] _04263_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ team_01_WB.instance_to_wrap.cpu.f0.state\[3\] _04505_ net564 vssd1 vssd1
+ vccd1 vccd1 _00019_ sky130_fd_sc_hd__a21o_1
X_15186_ net1180 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
X_12398_ net2510 net213 net426 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08775__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[41\] _04276_ _04295_ _04297_
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11349_ _05348_ _07224_ net346 _05347_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14068_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__nor2_1
XANTENNA__08527__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ net1165 team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] team_01_WB.instance_to_wrap.a1.WRITE_I
+ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21o_2
XANTENNA__12170__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17827_ clknet_leaf_88_wb_clk_i _03384_ _01648_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14886__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[30\] net720 _04800_
+ _04802_ _04810_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17758_ clknet_leaf_89_wb_clk_i net1824 _01579_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08884__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17472__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16709_ clknet_leaf_119_wb_clk_i _02269_ _00572_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_08491_ net999 net860 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and2_4
X_17689_ clknet_leaf_81_wb_clk_i _03249_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18197__1571 vssd1 vssd1 vccd1 vccd1 _18197__1571/HI net1571 sky130_fd_sc_hd__conb_1
XFILLER_0_45_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10357__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ _05364_ _05370_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ _05296_ _05301_ _05305_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__or4_4
XANTENNA__13339__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12345__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout309_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[27\] vssd1 vssd1 vccd1 vccd1
+ net2026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09558__A2 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__B team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold421 team_01_WB.instance_to_wrap.cpu.f0.num\[27\] vssd1 vssd1 vccd1 vccd1 net2037
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 net102 vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08766__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold454 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13965__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold465 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1120_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10092__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold476 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1218_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold498 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09945_ _06185_ _06192_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__nor3_2
XFILLER_0_25_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09881__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 _04670_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13176__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08518__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net947 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12080__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_4
X_09876_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__o21a_1
Xfanout967 _04501_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
Xhold1110 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] vssd1 vssd1 vccd1 vccd1
+ net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
Xhold1121 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[75\] vssd1 vssd1 vccd1 vccd1
+ net2748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\] net738 net701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a22o_1
XANTENNA__17815__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1176 team_01_WB.instance_to_wrap.cpu.K0.code\[5\] vssd1 vssd1 vccd1 vccd1 net2792
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net2803 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net1120 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] net913
+ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__and3_1
Xhold1198 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13814__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18081__1455 vssd1 vssd1 vccd1 vccd1 _18081__1455/HI net1455 sky130_fd_sc_hd__conb_1
XFILLER_0_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08689_ _04946_ _04948_ _04950_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__or4_1
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17965__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _06868_ _06981_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09121__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _05959_ _05923_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10267__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ team_01_WB.instance_to_wrap.cpu.f0.num\[28\] net328 net352 net1061 vssd1
+ vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10582_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] _04716_ vssd1 vssd1 vccd1
+ vccd1 _06846_ sky130_fd_sc_hd__nor2_1
XANTENNA__09797__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12321_ net3216 net264 net428 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12255__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net1251 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XANTENNA__11379__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net3236 net246 net435 vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__mux2_1
XANTENNA__08034__A team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ net511 _07403_ net529 vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__a21o_1
X_12183_ net2907 net279 net444 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__mux2_1
XANTENNA__10564__A0 _06826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ _06991_ _07171_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__nor2_1
XANTENNA__09791__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16991_ clknet_leaf_5_wb_clk_i _02551_ _00854_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11395__A _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15942_ net1342 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__inv_2
X_11065_ _05760_ _07199_ net324 vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__a21o_1
XANTENNA__10316__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] net883 vssd1
+ vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17495__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15873_ net1397 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__inv_2
XANTENNA__08367__A_N team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17612_ clknet_leaf_44_wb_clk_i _03172_ _01475_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14824_ net1350 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17543_ clknet_leaf_123_wb_clk_i _03103_ _01406_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14755_ net1183 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
X_11967_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__and2b_2
XANTENNA__13281__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13706_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] _04027_ vssd1 vssd1 vccd1 vccd1
+ _04028_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ net518 _07018_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__nand2_1
X_17474_ clknet_leaf_143_wb_clk_i _03034_ _01337_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14686_ net1378 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net3110 net210 net482 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13569__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16425_ clknet_leaf_86_wb_clk_i _02053_ _00288_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\]
+ sky130_fd_sc_hd__dfstp_1
X_13637_ _03805_ _03969_ _03804_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10849_ _05788_ _05852_ _05923_ _05993_ net506 net511 vssd1 vssd1 vccd1 vccd1 _07113_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14230__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16356_ clknet_leaf_66_wb_clk_i net1671 _00224_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13568_ net767 _07307_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09966__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15307_ net1210 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
X_12519_ net1958 net269 net410 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12165__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16287_ clknet_leaf_98_wb_clk_i _01921_ _00155_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ _03836_ _03840_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18026_ net1420 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ net1287 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XANTENNA__12544__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15169_ net1287 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10555__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08879__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout208 _07879_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
XFILLER_0_5_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16712__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 _07925_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
XFILLER_0_120_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09730_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] net668 vssd1 vssd1
+ vccd1 vccd1 _05994_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[11\] net887
+ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__and3_1
X_08612_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\] net736 net717 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09592_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\] net864 vssd1
+ vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09503__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08543_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\] net940 vssd1
+ vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_A _07989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08474_ net1108 net1111 net1114 net1106 vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10087__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__A1 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11035__B2 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16242__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17368__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10794__A0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1335_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] net950
+ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11338__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold240 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10546__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 _03398_ vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _01972_ vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold273 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\] vssd1 vssd1 vccd1 vccd1
+ net1889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold284 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1
+ net1900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout962_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout720 _04672_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_6
XFILLER_0_121_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout731 _04661_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_6
X_09928_ _06189_ _06190_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__or3_1
Xfanout742 net743 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout753 _04639_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_8
XFILLER_0_121_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout764 _04634_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
Xfanout786 _04511_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10849__A1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\] net926 vssd1
+ vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__and3_1
Xfanout797 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit vssd1 vssd1 vccd1 vccd1 net797
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13634__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15415__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ _03577_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08955__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13799__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11821_ _07855_ _07944_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13263__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ net1323 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XANTENNA__10077__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ net3118 net204 net481 vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10762__A_N net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10703_ net549 net521 net515 net501 vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__and4_1
X_14471_ net1335 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ team_01_WB.instance_to_wrap.cpu.K0.count\[0\] team_01_WB.instance_to_wrap.cpu.K0.enable
+ net1169 vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ clknet_leaf_117_wb_clk_i _01877_ _00078_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _03773_ _03774_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10634_ _06889_ _06895_ _06897_ _06891_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__a211o_1
X_17190_ clknet_leaf_139_wb_clk_i _02750_ _01053_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09786__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12774__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16141_ net1332 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08978__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13353_ net3 net801 net596 net2935 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a22o_1
X_10565_ _06807_ _06828_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__and2_1
XANTENNA__08442__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12304_ net3020 net202 net429 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__mux2_1
X_16072_ net1377 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__inv_2
X_13284_ net104 net815 net598 net1670 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16735__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10496_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\] net649 net639 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12526__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15023_ net1248 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
X_12235_ net2055 net192 net435 vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
XANTENNA__12713__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10537__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08699__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12166_ net3222 net213 net450 vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18196__1570 vssd1 vssd1 vccd1 vccd1 _18196__1570/HI net1570 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ _07380_ net324 _07346_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__or3b_1
XANTENNA__16885__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ net2300 net295 net458 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__mux2_1
X_16974_ clknet_leaf_50_wb_clk_i _02534_ _00837_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11048_ _07276_ _07280_ net522 vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__mux2_1
X_15925_ net1351 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__inv_2
XANTENNA__09026__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08902__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15325__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ net1253 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09323__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ net1380 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15787_ net1204 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__inv_2
XANTENNA__10469__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ net2929 net220 net362 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10068__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11265__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14738_ net1324 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
X_17526_ clknet_leaf_33_wb_clk_i _03086_ _01389_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08584__D net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17457_ clknet_leaf_20_wb_clk_i _03017_ _01320_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16265__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14669_ net1369 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08681__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16408_ clknet_leaf_103_wb_clk_i _02036_ _00271_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_08190_ _04584_ _04587_ _04589_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__or3_1
X_17388_ clknet_leaf_45_wb_clk_i _02948_ _01251_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08969__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16339_ clknet_leaf_64_wb_clk_i net1796 _00207_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09993__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18009_ clknet_leaf_84_wb_clk_i _03558_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12623__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18080__1454 vssd1 vssd1 vccd1 vccd1 _18080__1454/HI net1454 sky130_fd_sc_hd__conb_1
XANTENNA__14404__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10651__B _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09713_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] net930
+ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout376_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09644_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\] net743 _04656_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\] vssd1 vssd1 vccd1 vccd1
+ _05908_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17040__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09233__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ _05829_ _05836_ _05837_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1285_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] net643 _04789_
+ net672 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18025__1419 vssd1 vssd1 vccd1 vccd1 _18025__1419/HI net1419 sky130_fd_sc_hd__conb_1
X_08457_ net764 _04719_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__nor3_1
XFILLER_0_93_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08672__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08388_ net1147 net1151 net1153 net1149 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10767__A0 _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10350_ _06037_ _06605_ _05208_ _05488_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09009_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] net622 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10281_ net1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[0\] net866 vssd1
+ vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12533__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10842__A _06314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ net2261 net248 net463 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10280__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 net551 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14130__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13931__A_N net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_2
X_13971_ net1170 _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__nand2_2
Xfanout583 _04721_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_2
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_2
X_15710_ net1313 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
X_12922_ net2260 net604 net586 _03619_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a22o_1
X_16690_ clknet_leaf_55_wb_clk_i _02250_ _00553_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15641_ net1191 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11392__B _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12853_ net1924 net242 net368 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11804_ _07857_ _07930_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15572_ net1243 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
X_12784_ net2295 net263 net376 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08112__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17311_ clknet_leaf_5_wb_clk_i _02871_ _01174_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14523_ net1403 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
X_11735_ net2868 net193 net479 vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12708__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08663__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17242_ clknet_leaf_36_wb_clk_i _02802_ _01105_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14197__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14454_ net1392 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11666_ net1869 net1160 net568 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1
+ vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a22o_1
X_13405_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _06663_ vssd1 vssd1
+ vccd1 vccd1 _03758_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10617_ _06525_ _06880_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__nor2_1
X_17173_ clknet_leaf_25_wb_clk_i _02733_ _01036_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14385_ net1382 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
X_11597_ net496 _07813_ net2049 net838 vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16124_ net1395 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13336_ net21 net798 net593 net2704 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__o22a_1
X_10548_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] net646 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16055_ net1368 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13267_ net1842 net816 net600 team_01_WB.instance_to_wrap.a1.ADR_I\[24\] vssd1 vssd1
+ vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
XANTENNA__12443__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\] net739 net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15006_ net1300 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XANTENNA__09376__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ net2181 net275 net440 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12149_ net2732 net252 net449 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10930__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14121__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16957_ clknet_leaf_128_wb_clk_i _02517_ _00820_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10289__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ net1346 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16888_ clknet_leaf_26_wb_clk_i _02448_ _00751_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08595__C _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15839_ net1294 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__inv_2
XANTENNA__10199__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09988__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\] net930 vssd1
+ vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__and3_1
XANTENNA__08103__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10446__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11789__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[45\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
X_17509_ clknet_leaf_134_wb_clk_i _03069_ _01372_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_09291_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\] net955
+ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12618__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_13 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11841__A1_N net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08242_ net2283 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\] net1047 vssd1 vssd1
+ vccd1 vccd1 _03505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10646__B _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13022__B _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08173_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__or4b_2
XANTENNA__10749__A0 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10213__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12353__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_100_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__09906__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09228__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_A _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13184__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16430__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17556__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08342__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09627_ _05788_ _05822_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__nor2_1
XANTENNA__08893__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11229__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09558_ net581 _05820_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ net1003 net843 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__and2_4
XFILLER_0_13_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12528__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__A _06867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ _05719_ net558 net582 vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__mux2_2
XFILLER_0_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11520_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07713_ vssd1 vssd1 vccd1 vccd1
+ _07760_ sky130_fd_sc_hd__or2_1
XANTENNA__14179__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10452__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] team_01_WB.instance_to_wrap.cpu.f0.i\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10275__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire258 _07929_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_4
X_10402_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14170_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[99\] _04250_ _04276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\]
+ _04328_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11382_ _06776_ net339 _07492_ net542 _07645_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__a221oi_1
XANTENNA__09070__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13121_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\] net2387 net829 vssd1 vssd1
+ vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ _06385_ _06595_ _06384_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12263__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input54_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ net1678 _03687_ net1030 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
XANTENNA__09138__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[0\] net870 vssd1
+ vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__and3_1
XANTENNA__08042__A team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11165__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ net2911 net193 net463 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
Xfanout1301 net1302 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_4
X_10195_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[1\] net945 vssd1
+ vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__and3_1
X_17860_ clknet_leaf_78_wb_clk_i net1632 _01680_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1312 net1313 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__buf_4
Xfanout1323 net1325 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__buf_4
Xfanout1334 net1335 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__buf_4
XANTENNA__14103__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16811_ clknet_leaf_46_wb_clk_i _02371_ _00674_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1345 net1349 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__clkbuf_4
Xfanout1356 net1360 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__buf_2
X_17791_ clknet_leaf_70_wb_clk_i _03348_ _01612_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout1367 net1370 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1378 net1379 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__buf_4
Xfanout380 net382 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_6
Xfanout391 _03566_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_6
Xfanout1389 net1414 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13954_ _04509_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__nor2_1
X_16742_ clknet_leaf_141_wb_clk_i _02302_ _00605_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12905_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\] _07307_ net1032 vssd1 vssd1
+ vccd1 vccd1 _03607_ sky130_fd_sc_hd__mux2_1
X_16673_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[27\]
+ _00536_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13885_ _04124_ _04125_ team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\] _04144_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_atmax sky130_fd_sc_hd__and4_4
XANTENNA__11483__A4 _07734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15624_ net1209 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
X_12836_ net3067 net286 net367 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__mux2_1
XANTENNA__12968__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15555_ net1223 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XANTENNA__12968__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ net2022 net202 net377 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
XANTENNA__12438__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08636__A2 _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14506_ net1343 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
XANTENNA__10443__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11718_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _07858_ vssd1 vssd1
+ vccd1 vccd1 _07859_ sky130_fd_sc_hd__and2_1
X_15486_ net1300 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12698_ net3209 net190 net383 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__mux2_1
X_17225_ clknet_leaf_40_wb_clk_i _02785_ _01088_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14437_ net1387 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ net1743 net1157 net567 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1
+ vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a22o_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput44 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13393__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17156_ clknet_leaf_138_wb_clk_i _02716_ _01019_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14368_ net1326 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
Xinput55 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XANTENNA__16303__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput66 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_1
XANTENNA__17429__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold806 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ net1400 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold817 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ net135 net813 net807 net1784 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a22o_1
Xhold828 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\] vssd1 vssd1 vccd1 vccd1
+ net2455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12173__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17087_ clknet_leaf_1_wb_clk_i _02647_ _00950_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14299_ net1367 _04443_ _04444_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16038_ net1373 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__inv_2
XANTENNA_wire559_A _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16453__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08860_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\] net646 _05111_
+ _05118_ _05119_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10903__A0 _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18024__1418 vssd1 vssd1 vccd1 vccd1 _18024__1418/HI net1418 sky130_fd_sc_hd__conb_1
XFILLER_0_104_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1506 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net3122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net3133 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08791_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] net910 net640 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\]
+ net670 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__a221o_1
X_17989_ clknet_leaf_68_wb_clk_i _03538_ _01809_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1528 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1539 team_01_WB.instance_to_wrap.cpu.f0.num\[22\] vssd1 vssd1 vccd1 vccd1 net3155
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039__1429 vssd1 vssd1 vccd1 vccd1 _18039__1429/HI net1429 sky130_fd_sc_hd__conb_1
XANTENNA__08875__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] net652 _05657_
+ _05671_ _05672_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09343_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] net897
+ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12348__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08627__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A _07884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10434__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09274_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] net850 vssd1
+ vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18175__1549 vssd1 vssd1 vccd1 vccd1 _18175__1549/HI net1549 sky130_fd_sc_hd__conb_1
X_08225_ _04560_ _04618_ _04619_ net1036 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1150_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10095__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1248_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09588__B1 _05850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13384__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08156_ net1707 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1
+ vccd1 vccd1 _03539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09884__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12083__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] team_01_WB.instance_to_wrap.cpu.f0.num\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11147__B1 _07399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12811__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16946__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] net897
+ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09512__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10951_ _05551_ net335 net331 _05552_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09124__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08866__A2 _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13670_ net769 _03995_ net968 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a21oi_1
X_10882_ _06718_ net334 net332 _06719_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12621_ net2121 net316 net397 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13072__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__A _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15340_ net1263 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12552_ net1910 net267 net406 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08037__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _07743_ _07748_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15271_ net1182 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
X_12483_ net3233 net274 net412 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17010_ clknet_leaf_39_wb_clk_i _02570_ _00873_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09579__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14222_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\] _04249_ _04252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\]
+ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a221o_1
XANTENNA__13375__B2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] _07689_ vssd1 vssd1 vccd1
+ vccd1 _07692_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14153_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] _04253_ _04268_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[42\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a22o_1
XANTENNA__16476__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11365_ _07070_ _07076_ _07336_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13104_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[4\] _06313_ net1036 vssd1
+ vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10316_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] net696 net688 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14084_ _04226_ net789 _04243_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__and3_4
XFILLER_0_24_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output160_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ _06998_ _07475_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__or2_1
X_13035_ net2631 net834 net354 _03676_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a22o_1
X_17912_ clknet_leaf_101_wb_clk_i net2940 _01732_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] net618 _06496_ _06501_
+ _06503_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12721__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1120 net1123 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1131 net1133 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09751__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17843_ clknet_leaf_80_wb_clk_i net1940 _01663_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1142 net1146 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_4
X_10178_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] net615 _06425_ _06426_
+ _06439_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08500__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1153 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1 vccd1
+ net1153 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17871__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1164 net1168 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1175 net1176 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_2
Xfanout1186 net1194 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_4
X_17774_ clknet_leaf_105_wb_clk_i _03332_ _01595_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1197 net1203 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_4
XFILLER_0_135_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10327__A1_N net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14986_ net1202 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16725_ clknet_leaf_26_wb_clk_i _02285_ _00588_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13937_ net1164 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[18\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[18\] sky130_fd_sc_hd__and3b_1
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17101__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13868_ _04506_ team_01_WB.instance_to_wrap.a1.READ_I team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ _04508_ team_01_WB.instance_to_wrap.a1.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _00009_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16656_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[10\]
+ _00519_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09331__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11580__B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ net2474 net314 net372 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__mux2_1
X_15607_ net1239 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12168__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ net563 _07774_ _04100_ net786 vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16587_ clknet_leaf_89_wb_clk_i _02215_ _00450_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13602__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11613__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15538_ net1175 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09282__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15469_ net1213 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17208_ clknet_leaf_29_wb_clk_i _02768_ _01071_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09034__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18188_ net1562 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
XFILLER_0_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold603 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17139_ clknet_leaf_21_wb_clk_i _02699_ _01002_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 net2252
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09961_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\] net893 vssd1
+ vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold669 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08912_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\] net894
+ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09892_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\] net852 vssd1
+ vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__and3_1
XANTENNA__12877__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12631__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14412__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09506__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\] net885 vssd1
+ vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__and3_1
Xhold1303 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08410__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A _07874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1314 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1336 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2952 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout289_A _07901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1347 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
X_08774_ _05020_ _05035_ _05036_ _05037_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or4_1
Xhold1358 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11771__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12078__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout623_A _04768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1365_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\] net860
+ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16499__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] net885
+ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12806__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17744__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13357__A1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08208_ _04565_ _04573_ _04584_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__or4b_2
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09188_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] net842 vssd1
+ vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08139_ team_01_WB.instance_to_wrap.cpu.K0.keyvalid _04565_ vssd1 vssd1 vccd1 vccd1
+ _04566_ sky130_fd_sc_hd__and2_2
XFILLER_0_121_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11150_ _06870_ _07412_ _07413_ _07411_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__o211a_1
XANTENNA__10591__A1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\] net645 _04755_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a22o_1
XANTENNA__10591__B2 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11081_ _06888_ _06894_ _06600_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12541__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] net880 vssd1
+ vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__and3_1
XANTENNA__10343__A1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17124__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ net1341 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net1243 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
X_11983_ net2174 net251 net468 vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
X_13722_ _04021_ _04040_ _04558_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21oi_1
X_16510_ clknet_leaf_80_wb_clk_i net2209 _00373_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10934_ _06899_ _06900_ _06914_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__a21o_1
XANTENNA__11843__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17490_ clknet_leaf_39_wb_clk_i _03050_ _01353_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09789__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17274__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16441_ clknet_leaf_99_wb_clk_i _02069_ _00304_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[53\]
+ sky130_fd_sc_hd__dfstp_1
X_13653_ _03793_ _03809_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__xor2_1
XANTENNA__10297__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10865_ _06722_ _07128_ net322 vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12604_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\] net232 net396 vssd1
+ vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
XANTENNA__13596__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16372_ clknet_leaf_113_wb_clk_i net1619 _00240_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13584_ _03834_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and2_1
XANTENNA__08990__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10796_ net520 net514 _07058_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18023__1417 vssd1 vssd1 vccd1 vccd1 _18023__1417/HI net1417 sky130_fd_sc_hd__conb_1
X_15323_ net1316 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18111_ net1485 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12535_ net2950 net240 net405 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12716__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18042_ net1604 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_15254_ net1258 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12466_ net1960 net194 net413 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14205_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\] _04229_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\]
+ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11417_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _07679_ _07675_ vssd1
+ vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__mux2_1
X_15185_ net1196 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
X_12397_ net2278 net291 net424 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
XANTENNA__10463__C _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18038__1428 vssd1 vssd1 vccd1 vccd1 _18038__1428/HI net1428 sky130_fd_sc_hd__conb_1
X_14136_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\] _04268_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\]
+ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _06924_ _07228_ net323 vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15328__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12451__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ net792 net791 net790 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__and3_4
XFILLER_0_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11279_ _06997_ _07173_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13018_ net3103 net211 net363 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__mux2_1
XANTENNA__09326__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18174__1548 vssd1 vssd1 vccd1 vccd1 _18174__1548/HI net1548 sky130_fd_sc_hd__conb_1
X_17826_ clknet_leaf_79_wb_clk_i _03383_ _01647_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17757_ clknet_leaf_115_wb_clk_i _03315_ _01578_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ net1192 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15063__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16708_ clknet_leaf_129_wb_clk_i _02268_ _00571_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08490_ net1107 net1109 net1112 net1115 vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__and4_4
X_17688_ clknet_leaf_76_wb_clk_i _03248_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15998__A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[25\]
+ _00502_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17767__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09996__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09111_ _05371_ _05372_ _05373_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08463__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09042_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] net741 net727 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\]
+ _05291_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a221o_1
XANTENNA__09007__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08405__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16791__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout204_A _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\] vssd1 vssd1 vccd1 vccd1
+ net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold455 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17147__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ _06196_ _06199_ _06203_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__or4_1
Xhold488 net148 vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold499 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1 vccd1
+ net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net915 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 net926 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_4
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_2
X_09875_ net713 _06129_ _06134_ _06138_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__or4_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 net959 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_4
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_2
Xhold1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A _07803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1111 _03449_ vssd1 vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net993 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_2
Xhold1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\] net749 _05073_
+ _05077_ _05079_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a2111o_1
Xhold1133 _02099_ vssd1 vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10876__A2 _07139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16171__CLK clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1155 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17297__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1177 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] net920 vssd1
+ vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13275__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1188 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13192__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout838_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08688_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] net657 net630 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\]
+ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09402__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10650_ _06043_ _06912_ _06913_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09309_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] net751 net712 _05560_
+ _05563_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12536__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net1155 _06844_ vssd1 vssd1 vccd1
+ vccd1 _06845_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[11\] net267 net429 vssd1
+ vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08206__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net1961 net277 net437 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10013__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ net517 _07434_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ net2445 net250 net445 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11133_ _06600_ _06888_ _06894_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12271__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16990_ clknet_leaf_4_wb_clk_i _02550_ _00853_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13502__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16514__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ net1340 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11064_ _05760_ _07199_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__nor2_1
XANTENNA__08050__A team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ net581 _06278_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__or2_1
X_15872_ net1397 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17611_ clknet_leaf_60_wb_clk_i _03171_ _01474_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14823_ net1354 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XANTENNA__13266__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13805__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16664__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17542_ clknet_leaf_139_wb_clk_i _03102_ _01405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14754_ net1274 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
X_11966_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__and2_2
XANTENNA__09485__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13705_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _04026_ vssd1 vssd1 vccd1 vccd1
+ _04027_ sky130_fd_sc_hd__or2_1
X_10917_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17473_ clknet_leaf_136_wb_clk_i _03033_ _01336_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14685_ net1375 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11897_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _04622_ _08005_ _08006_
+ vssd1 vssd1 vccd1 vccd1 _08007_ sky130_fd_sc_hd__a22o_1
XANTENNA__14215__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13569__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16424_ clknet_leaf_105_wb_clk_i _02052_ _00287_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\]
+ sky130_fd_sc_hd__dfstp_1
X_13636_ _03793_ _03809_ _03807_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10848_ net523 _07108_ net535 vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09237__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14230__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16355_ clknet_leaf_75_wb_clk_i net1624 _00223_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12446__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ _07908_ _03910_ net186 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ _07033_ _07042_ net538 vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12518_ net1844 net272 net407 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
X_15306_ net1201 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16286_ clknet_leaf_98_wb_clk_i _01920_ _00154_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13498_ _03846_ _03849_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18025_ net1419 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15237_ net1229 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
X_12449_ net1941 net217 net415 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10193__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15168_ net1273 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10555__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14119_ net792 _04237_ _04243_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__and3_4
XANTENNA__12181__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15099_ net1317 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
Xfanout209 _07879_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_1
XFILLER_0_10_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16194__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10921__C _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08598__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ _04719_ _04720_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1
+ vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09490__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08611_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\] _04676_ net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a22o_1
X_17809_ clknet_leaf_69_wb_clk_i _03366_ _01630_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09591_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\] net868 vssd1
+ vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08542_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\] net936
+ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10649__B _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08473_ net1018 net898 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08684__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10491__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14221__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11035__A2 _07033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12356__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout321_A _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10794__A1 _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] net941
+ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1230_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold230 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net1846
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 net123 vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[2\] vssd1 vssd1 vccd1 vccd1
+ net1868 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09892__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold263 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold274 _02136_ vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12091__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold285 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _04679_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_2
Xfanout721 _04671_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_8
Xfanout732 _04661_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09927_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\] net728 net726 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout743 _04651_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_8
XFILLER_0_42_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout754 _04639_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_2
X_18022__1416 vssd1 vssd1 vccd1 vccd1 _18022__1416/HI net1416 sky130_fd_sc_hd__conb_1
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_2
X_09858_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\] net941 vssd1
+ vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__and3_1
Xfanout787 _04231_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_2
XANTENNA__10849__A2 _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 net800 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
X_08809_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] net956
+ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and3_1
X_09789_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] net914 vssd1
+ vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11820_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _07854_ vssd1 vssd1
+ vccd1 vccd1 _07944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18037__1427 vssd1 vssd1 vccd1 vccd1 _18037__1427/HI net1427 sky130_fd_sc_hd__conb_1
X_11751_ net774 _07885_ _07886_ _07887_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__08675__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13650__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ net549 net500 vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14470_ net1336 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11682_ net1169 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.next_state
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14212__A2 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13421_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net591 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__a21o_1
X_10633_ _06178_ _06896_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17312__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ net1314 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13352_ net4 net798 net593 net3190 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__o22a_1
X_10564_ _06826_ _06827_ net578 vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__mux2_1
X_18173__1547 vssd1 vssd1 vccd1 vccd1 _18173__1547/HI net1547 sky130_fd_sc_hd__conb_1
XANTENNA__08045__A team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ net2179 net240 net429 vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XANTENNA__13886__A team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16071_ net1368 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13283_ net105 net813 net599 net1642 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10495_ _06757_ _06758_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__or2_1
X_15022_ net1231 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XANTENNA__09927__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ net2152 net194 net436 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
XANTENNA__17462__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12165_ net2394 net291 net448 vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ _06179_ _06892_ _07345_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12096_ net2846 net309 net458 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__mux2_1
X_16973_ clknet_leaf_21_wb_clk_i _02533_ _00836_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11047_ net532 _07097_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nand2_1
X_15924_ net1351 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13239__A0 _03723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__B2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15855_ net1248 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ net1343 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
X_15786_ net1199 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__inv_2
X_12998_ net3200 net283 net360 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17525_ clknet_leaf_26_wb_clk_i _03085_ _01388_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14737_ net1323 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
X_11949_ net2590 net278 net472 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15341__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17456_ clknet_leaf_24_wb_clk_i _03016_ _01319_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14668_ net1373 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14203__A2 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08881__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ clknet_leaf_75_wb_clk_i _02035_ _00270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12176__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ _03815_ _03947_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__nor2_1
X_17387_ clknet_leaf_51_wb_clk_i _02947_ _01250_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ net1371 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16338_ clknet_leaf_62_wb_clk_i net1878 _00206_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17805__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16269_ clknet_leaf_69_wb_clk_i _01906_ _00137_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ clknet_leaf_84_wb_clk_i _03557_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09918__B1 _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09712_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] net940
+ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09643_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\] net915 vssd1
+ vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout271_A _07957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout369_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] net720 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\]
+ _05825_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__a221o_1
XANTENNA__09449__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08525_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[31\] net641 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout536_A _06383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10098__C net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17335__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1278_A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08456_ _04487_ net765 net682 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a21o_2
XFILLER_0_110_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09887__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ net1117 net948 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and2_4
XANTENNA__12086__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10216__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17485__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A1 _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12814__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _05268_ _05269_ _05270_ _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__or4_1
X_10280_ net1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] net899 vssd1
+ vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09127__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _06382_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_2
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_2
XANTENNA__15426__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ net584 vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__mux2_1
Xfanout573 _07803_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_2
Xfanout584 _04157_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout595 _03748_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
XANTENNA__09424__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] net1053 net364 _03618_
+ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08896__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15640_ net1255 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
X_12852_ net2539 net316 net368 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _07856_ vssd1 vssd1
+ vccd1 vccd1 _07930_ sky130_fd_sc_hd__nor2_1
X_12783_ net2185 net269 net378 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
X_15571_ net1179 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11247__A2 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12444__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17310_ clknet_leaf_3_wb_clk_i _02870_ _01173_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14522_ net1407 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11734_ net774 _07871_ _07873_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16702__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17241_ clknet_leaf_17_wb_clk_i _02801_ _01104_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14453_ net1392 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
X_11665_ net1690 net1160 net568 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1
+ vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10207__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10616_ net505 _06591_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__nor2_1
X_13404_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] _04955_ vssd1 vssd1
+ vccd1 vccd1 _03757_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14384_ net1329 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
X_17172_ clknet_leaf_9_wb_clk_i _02732_ _01035_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[28\] net572 vssd1 vssd1 vccd1
+ vccd1 _07813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16123_ net1395 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__inv_2
X_13335_ net22 net798 net593 net2669 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10547_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\] net653 net628 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\]
+ _06810_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__a221o_1
XANTENNA__12724__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17978__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13266_ net92 net816 net600 net1620 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
X_16054_ net1373 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__inv_2
X_10478_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] net754 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\]
+ _06728_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__a221o_1
XANTENNA__08503__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15005_ net1282 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
X_12217_ net2328 net216 net439 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13197_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[45\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__C net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ net3088 net255 net448 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net2006 net282 net455 vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
X_16956_ clknet_leaf_15_wb_clk_i _02516_ _00819_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08876__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ net1345 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08887__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16887_ clknet_leaf_12_wb_clk_i _02447_ _00750_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16232__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11075__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15838_ net1315 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15769_ net1191 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
X_08310_ net2508 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\] net1041 vssd1 vssd1
+ vccd1 vccd1 _03437_ sky130_fd_sc_hd__mux2_1
X_17508_ clknet_leaf_128_wb_clk_i _03068_ _01371_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_09290_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\] net953 vssd1
+ vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08241_ net2352 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03506_ sky130_fd_sc_hd__mux2_1
XANTENNA_14 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ clknet_leaf_4_wb_clk_i _02999_ _01302_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09500__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08172_ _04551_ _04570_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10749__A1 _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12634__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14415__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__S1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_100_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1026_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13871__B1 _04617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A _04743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18172__1546 vssd1 vssd1 vccd1 vccd1 _18172__1546/HI net1546 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1395_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ _05852_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__nand2_2
XFILLER_0_74_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net591 net581 vssd1 vssd1
+ vccd1 vccd1 _05821_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout820_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12809__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10437__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ net1107 net1115 net1112 net1109 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09488_ net558 vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__inv_2
XANTENNA__10837__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08439_ _04700_ _04701_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16875__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\] team_01_WB.instance_to_wrap.cpu.f0.i\[29\]
+ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10401_ _06643_ _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nand2_1
XANTENNA__12544__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11381_ _06778_ net342 net334 _06774_ _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10853__A _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13120_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\] net2208 net827 vssd1 vssd1
+ vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10332_ _06385_ _06595_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _05063_ net571 net359 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__o21a_1
X_10263_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] net862 vssd1
+ vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10291__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ net2251 net196 net465 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__mux2_1
Xfanout1302 net1415 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input47_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\] net932 vssd1
+ vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1313 net1314 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__clkbuf_4
Xfanout1324 net1325 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16255__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__B2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16810_ clknet_leaf_43_wb_clk_i _02370_ _00673_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1335 net1337 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__buf_4
XANTENNA__08581__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1346 net1348 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__buf_4
X_17790_ clknet_leaf_116_wb_clk_i net1157 _01611_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.pc_enable
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1357 net1359 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__buf_4
Xfanout370 _03572_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_4
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1368 net1370 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__buf_4
XANTENNA__08696__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1379 net1414 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__buf_2
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_4
Xfanout392 _03566_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_4
X_16741_ clknet_leaf_134_wb_clk_i _02301_ _00604_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13953_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _04146_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12904_ net1618 net607 net589 _03606_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16672_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[26\]
+ _00535_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ team_01_WB.instance_to_wrap.cpu.c0.count\[3\] team_01_WB.instance_to_wrap.cpu.c0.count\[2\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.next_count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__A2 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17650__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15623_ net1195 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
X_12835_ net3069 net231 net367 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12719__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08097__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13404__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15554_ net1286 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
X_12766_ net2730 net240 net377 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09833__A2 _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505_ net1343 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
X_11717_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__and3_1
X_15485_ net1283 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
X_12697_ net3031 net194 net385 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
XANTENNA__10466__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17224_ clknet_leaf_45_wb_clk_i _02784_ _01087_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14436_ net1212 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
X_11648_ net1159 _07835_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__nor2_1
XANTENNA__12962__B _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput45 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17155_ clknet_leaf_119_wb_clk_i _02715_ _01018_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11579_ _07731_ _07796_ _07801_ _07700_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__a32o_1
XANTENNA__12454__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14367_ net1326 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
Xinput56 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
Xinput67 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xhold807 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ net1388 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__inv_2
Xhold818 team_01_WB.instance_to_wrap.cpu.c0.count\[11\] vssd1 vssd1 vccd1 vccd1 net2434
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09329__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13318_ net136 net814 net807 net1701 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a22o_1
X_14298_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\]
+ _04195_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17086_ clknet_leaf_3_wb_clk_i _02646_ _00949_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16037_ net1355 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__inv_2
X_13249_ net47 net49 net48 net46 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__or4b_2
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18119__1493 vssd1 vssd1 vccd1 vccd1 _18119__1493/HI net1493 sky130_fd_sc_hd__conb_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09990__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10903__A1 _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08572__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1507 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3123 sky130_fd_sc_hd__dlygate4sd3_1
X_08790_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[22\] net658 net624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a22o_1
X_17988_ clknet_leaf_56_wb_clk_i _03537_ _01808_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1518 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net3134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 team_01_WB.instance_to_wrap.a1.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1 net3145
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16748__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16939_ clknet_leaf_46_wb_clk_i _02499_ _00802_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09411_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[13\] net642 net625 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12629__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09342_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] net845
+ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10419__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08408__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11092__A0 _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] net882
+ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__and3_1
XANTENNA__09230__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11631__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08224_ team_01_WB.instance_to_wrap.cpu.f0.state\[2\] team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13968__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09588__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08155_ net1807 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1
+ vccd1 vccd1 _03540_ sky130_fd_sc_hd__a22o_1
XANTENNA__11769__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1143_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ team_01_WB.instance_to_wrap.cpu.f0.i\[31\] team_01_WB.instance_to_wrap.cpu.f0.num\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17523__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1310_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1408_A net1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout868_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14097__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net1084 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[19\] net872
+ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__and3_1
XANTENNA__17673__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09405__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15704__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _06992_ _06999_ _07107_ _07212_ _07213_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__a32o_1
XANTENNA__10122__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09702__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09609_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\] net904 vssd1
+ vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10881_ _07143_ _07144_ _07142_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12539__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__A2_N net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12620_ net2798 net305 net398 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12551_ net1959 net270 net403 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11502_ net1062 _07720_ _07745_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1
+ vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__a31o_1
XANTENNA__10286__C _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15270_ net1281 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12482_ net2433 net215 net411 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11433_ _07691_ net1826 _07685_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__mux2_1
X_14221_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\] _04238_ _04260_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\]
+ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a22o_1
XANTENNA__12274__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\] _04255_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__a22o_1
X_11364_ _06942_ _07627_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08053__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ net1784 net837 net357 _03721_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[0\] net737 _06562_ _06566_
+ _06572_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__a2111o_1
X_14083_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] _04242_ _04244_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\]
+ _04240_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _06954_ _07555_ _07558_ _07106_ _07557_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__a221oi_1
XANTENNA__11138__A1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13034_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\] _03675_ net1028 vssd1
+ vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__mux2_1
X_17911_ clknet_leaf_108_wb_clk_i _03461_ _01731_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_10246_ _06493_ _06494_ _06498_ _06500_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12886__B2 _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[22\] vssd1 vssd1 vccd1 vccd1
+ net1110 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08554__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__A0 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_2
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_2
X_17842_ clknet_leaf_79_wb_clk_i net2299 _01662_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10177_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\] net649 _06423_ _06424_
+ _06429_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__a2111o_1
Xfanout1143 net1146 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08500__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1154 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1 vccd1
+ net1154 sky130_fd_sc_hd__buf_1
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_2
Xfanout1176 net1185 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
X_17773_ clknet_leaf_95_wb_clk_i _03331_ _01594_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14985_ net1210 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
Xfanout1187 net1194 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
Xfanout1198 net1203 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15614__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724_ clknet_leaf_4_wb_clk_i _02284_ _00587_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13936_ net1168 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[17\] sky130_fd_sc_hd__and3b_1
XFILLER_0_92_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09612__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__B _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16655_ clknet_leaf_96_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[9\]
+ _00518_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13867_ team_01_WB.instance_to_wrap.a1.WRITE_I _04507_ team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ _04508_ net2658 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a32o_1
XANTENNA__12449__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ net1304 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
XANTENNA__13063__A1 _05344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12818_ net3060 net302 net371 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
X_16586_ clknet_leaf_72_wb_clk_i _02214_ _00449_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13798_ _04475_ _07772_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13944__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14260__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15537_ net1196 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09050__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12749_ net3109 net270 net379 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
XANTENNA__12973__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10196__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15468_ net1262 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XANTENNA__09985__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17207_ clknet_leaf_10_wb_clk_i _02767_ _01070_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14419_ net1279 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18187_ net1561 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
XANTENNA__12184__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15399_ net1182 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18171__1545 vssd1 vssd1 vccd1 vccd1 _18171__1545/HI net1545 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17138_ clknet_leaf_31_wb_clk_i _02698_ _01001_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold604 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\] vssd1 vssd1 vccd1 vccd1
+ net2220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold637 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ clknet_leaf_53_wb_clk_i _02629_ _00932_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_09960_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] net848 vssd1
+ vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__and3_1
Xhold659 team_01_WB.instance_to_wrap.a1.ADR_I\[31\] vssd1 vssd1 vccd1 vccd1 net2275
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\] net849
+ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__and3_1
X_09891_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\] net879 vssd1
+ vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and3_1
XANTENNA__12877__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08842_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] net893
+ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__and3_1
Xhold1304 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08410__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1315 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1326 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08773_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\] net724 net720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__a22o_1
Xhold1337 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09225__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1359 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12359__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1093_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout449_A _08019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13054__A1 _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14251__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\] net909
+ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11065__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12883__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1260_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] net885 vssd1
+ vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09895__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08207_ _04553_ _04571_ _04572_ _04564_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13357__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ net1078 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\] net867
+ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__and3_1
XANTENNA__12094__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11368__A1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _04551_ _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16913__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13109__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__A1 _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ team_01_WB.instance_to_wrap.cpu.f0.num\[2\] vssd1 vssd1 vccd1 vccd1 _04500_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12822__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10100_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\] net862 vssd1
+ vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap890 _04742_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_2
X_11080_ _07325_ _07327_ _07343_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__o21a_2
XFILLER_0_80_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08601__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\] net862 vssd1
+ vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_1676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16240__D _00020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10343__A2 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09135__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14770_ net1303 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ net2926 net256 net467 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
XANTENNA__08747__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ team_01_WB.instance_to_wrap.cpu.f0.i\[26\] _04020_ vssd1 vssd1 vccd1 vccd1
+ _04040_ sky130_fd_sc_hd__nand2_1
XANTENNA__09432__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10933_ net344 _07156_ _07195_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12269__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ clknet_leaf_106_wb_clk_i _02068_ _00303_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__13045__A1 _06826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ _06778_ _07126_ _06938_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__o21ai_1
X_13652_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] _03982_ net1067 vssd1
+ vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08048__A team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12603_ net2566 net236 net395 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16371_ clknet_leaf_76_wb_clk_i _02005_ _00239_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18118__1492 vssd1 vssd1 vccd1 vccd1 _18118__1492/HI net1492 sky130_fd_sc_hd__conb_1
XANTENNA__13596__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ net516 _07058_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__nand2_1
X_13583_ _03829_ _03838_ _03831_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__o21a_1
XANTENNA__16443__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18110_ net1484 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__11901__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15322_ net1303 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ net3041 net208 net405 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13348__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18041_ net1603 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_83_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15253_ net1177 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12465_ _07841_ _07846_ net489 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14204_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\] _04239_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__a22o_1
XANTENNA__11202__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ net769 _07121_ net187 _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__a2bb2o_1
X_12396_ net2120 net297 net426 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15184_ net1262 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
X_14135_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[57\] _04244_ _04275_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\]
+ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11347_ _07602_ _07604_ _07610_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08775__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12732__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09607__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14066_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__and2b_1
X_11278_ _05758_ net341 net331 _05689_ _07541_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__o221a_1
XANTENNA__08511__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] net871 vssd1
+ vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__and3_1
X_13017_ net3153 net290 net362 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11531__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11531__B2 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17825_ clknet_leaf_80_wb_clk_i _03382_ _01646_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1 team_01_WB.instance_to_wrap.cpu.K0.state vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11872__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17756_ clknet_leaf_115_wb_clk_i _03314_ _01577_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.bit30
+ sky130_fd_sc_hd__dfrtp_4
X_14968_ net1254 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
XANTENNA__13284__B2 net1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09342__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16707_ clknet_leaf_119_wb_clk_i _02267_ _00570_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08884__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13919_ net1165 net1059 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[0\] sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17687_ clknet_leaf_84_wb_clk_i _03247_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11834__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12179__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ net1190 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XANTENNA__13036__A1 _06662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16638_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[24\]
+ _00501_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14233__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16569_ clknet_leaf_126_wb_clk_i _02197_ _00432_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09110_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\] net716 _05353_ _05354_
+ _05360_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09660__B1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16936__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09041_ _05302_ _05303_ _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__or3_1
X_18239_ net601 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13339__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08405__B net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold401 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold412 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold423 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 team_01_WB.instance_to_wrap.cpu.c0.count\[2\] vssd1 vssd1 vccd1 vccd1 net2050
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[48\] vssd1 vssd1 vccd1 vccd1
+ net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12642__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold456 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold467 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[23\] vssd1 vssd1 vccd1 vccd1
+ net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold489 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] net723 _06204_ _06205_
+ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08421__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_4
XANTENNA__08518__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09874_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\] _04656_ _06135_
+ _06136_ _06137_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a2111o_1
Xfanout947 _04652_ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_4
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
Xhold1101 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 _04501_ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
Xhold1112 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\] net719 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\]
+ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a221o_1
Xhold1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _04202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\] vssd1 vssd1 vccd1 vccd1
+ net2761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11782__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1178 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] net746 net701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a22o_1
XANTENNA__13275__B2 team_01_WB.instance_to_wrap.a1.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[58\] vssd1 vssd1 vccd1 vccd1
+ net2805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09252__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12089__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\] _04759_ net611
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[28\] vssd1 vssd1 vccd1 vccd1
+ _04951_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout733_A _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13027__A1 _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14224__B1 _04246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12817__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09308_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\] net725 net715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\]
+ _05558_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _04486_ vssd1 vssd1 vccd1
+ vccd1 _06844_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17861__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09239_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\] net745 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\]
+ _05497_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12250_ net1930 net217 net435 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ _07206_ _07360_ net522 vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__mux2_1
X_12181_ net2048 net255 net444 vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__mux2_1
XANTENNA__12552__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A1 _07653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ net345 _07349_ _07395_ _07394_ _07381_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__o311a_2
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09427__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15940_ net1340 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ net346 _07326_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10316__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] net765 _04723_ net1098 vssd1
+ vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__a22o_1
X_15871_ net1397 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__inv_2
X_17610_ clknet_leaf_41_wb_clk_i _03170_ _01473_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16809__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14822_ net1354 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09162__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17541_ clknet_leaf_129_wb_clk_i _03101_ _01404_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11277__B1 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18170__1544 vssd1 vssd1 vccd1 vccd1 _18170__1544/HI net1544 sky130_fd_sc_hd__conb_1
X_14753_ net1228 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11965_ net3251 net213 net474 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17391__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13704_ _04464_ _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17472_ clknet_leaf_142_wb_clk_i _03032_ _01335_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _07012_ _07016_ net512 vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14215__B1 _04372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14684_ net1399 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
X_11896_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\] net677 net779 vssd1 vssd1
+ vccd1 vccd1 _08006_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16959__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16423_ clknet_leaf_77_wb_clk_i _02051_ _00286_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_13635_ net969 _03968_ _03964_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12727__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10847_ net511 _07037_ _07100_ _07110_ net523 vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__o311a_1
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16354_ clknet_leaf_85_wb_clk_i _01988_ _00222_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ _03845_ _03903_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ _07036_ _07041_ net530 vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15305_ net1206 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12517_ net2051 net247 net409 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16285_ clknet_leaf_98_wb_clk_i _01919_ _00153_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13497_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _05134_ vssd1 vssd1
+ vccd1 vccd1 _03850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18024_ net1418 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15236_ net1269 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
X_12448_ net1856 net280 net416 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15167_ net1294 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
XANTENNA__12462__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ net2639 net219 net423 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
XANTENNA__09337__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ net792 net787 _04237_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__and3_4
X_15098_ net1258 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14049_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] _04215_ net566 vssd1
+ vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09173__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[29\] net732 net727 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a22o_1
X_17808_ clknet_leaf_68_wb_clk_i _03365_ _01629_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09590_ net580 _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\] net924
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__and3_1
X_17739_ clknet_leaf_96_wb_clk_i _03297_ _01560_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09503__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ net1106 net1109 net1115 net1112 vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__nor4b_1
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14206__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17884__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12637__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08416__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17114__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09024_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\] net949 vssd1
+ vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1056_A team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_01_WB.instance_to_wrap.a1.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net1836
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 net1847
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold242 _01974_ vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10546__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1223_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold253 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\] vssd1 vssd1 vccd1 vccd1
+ net1869 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12940__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold264 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17264__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout683_A _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold286 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\] vssd1 vssd1 vccd1 vccd1
+ net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _04685_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_6
Xhold297 team_01_WB.instance_to_wrap.a1.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1 net1913
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout711 net714 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_8
X_09926_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\] _04646_ _04656_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] vssd1 vssd1 vccd1 vccd1
+ _06190_ sky130_fd_sc_hd__a22o_1
Xfanout722 _04671_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout733 _04660_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_6
Xfanout744 _04648_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_8
X_18117__1491 vssd1 vssd1 vccd1 vccd1 _18117__1491/HI net1491 sky130_fd_sc_hd__conb_1
Xfanout755 net758 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_2
Xfanout766 _04630_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_2
X_09857_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\] net958 vssd1
+ vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__and3_1
Xfanout777 _04623_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_2
XANTENNA_fanout850_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 _04230_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_2
XANTENNA__10849__A3 _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout948_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ net976 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] net921 vssd1
+ vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__and3_1
X_09788_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\] net942 vssd1
+ vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08739_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[23\] net658 net640 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] net674 net774 vssd1 vssd1
+ vccd1 vccd1 _07887_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09872__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09710__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10701_ _04935_ _04883_ net501 vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__mux2_1
X_11681_ net37 net36 net35 net34 vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__nor4_2
XANTENNA__12547__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14328__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13420_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ net591 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _06175_ _06141_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ net1098 net763 net590 vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ net5 net798 net593 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1
+ vccd1 vccd1 _01929_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ net2814 net207 net429 vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16070_ net1374 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ net1997 net814 net599 net1829 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a22o_1
X_10494_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\] net643 net615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\]
+ _06755_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ net1213 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12282__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ _07842_ net494 _08011_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__and3_4
XANTENNA__10537__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12164_ net3242 net295 net450 vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
XANTENNA__09157__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08699__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11115_ net346 _07369_ _07370_ _07372_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__a311o_2
XFILLER_0_97_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ net3071 net312 net457 vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
X_16972_ clknet_leaf_44_wb_clk_i _02532_ _00835_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16631__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08996__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13487__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11046_ net322 _07126_ _07309_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__and3b_1
XFILLER_0_21_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15923_ net1360 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__inv_2
XANTENNA__11498__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15854_ net1230 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14805_ net1344 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XANTENNA__09323__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15785_ net1206 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12997_ net2471 net224 net361 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XANTENNA__10469__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17524_ clknet_leaf_6_wb_clk_i _03084_ _01387_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14736_ net1323 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
X_11948_ net2340 net252 net473 vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11670__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17455_ clknet_leaf_18_wb_clk_i _03015_ _01318_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12457__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14667_ net1363 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11879_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\] _07426_ net677 vssd1 vssd1
+ vccd1 vccd1 _07993_ sky130_fd_sc_hd__mux2_1
X_16406_ clknet_leaf_83_wb_clk_i net2280 _00269_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13618_ net969 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1
+ vccd1 _03954_ sky130_fd_sc_hd__nand2_1
X_17386_ clknet_leaf_42_wb_clk_i _02946_ _01249_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14598_ net1378 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16337_ clknet_leaf_63_wb_clk_i net1972 _00205_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08969__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13549_ net767 _07653_ net1066 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11973__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16161__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16268_ clknet_leaf_66_wb_clk_i _01905_ _00136_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09993__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18007_ clknet_leaf_84_wb_clk_i _03556_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15069__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15219_ net1186 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12192__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16199_ clknet_leaf_97_wb_clk_i _01866_ _00067_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12922__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12920__S net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09711_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[10\] net913
+ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__and3_1
XANTENNA__09146__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] net918
+ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09573_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] net748 net702 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__a22o_1
XANTENNA__09233__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08524_ _04781_ _04783_ _04785_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__or4_1
XANTENNA__12984__A1_N _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09530__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12367__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11661__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ net772 _04715_ net681 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout431_A _08023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout529_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08386_ net1151 net1153 net1147 net1149 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__and4b_4
XANTENNA__16504__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1340_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout898_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\] net656 _05246_
+ _05250_ _05255_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_108_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16654__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09408__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12830__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13469__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout530 _06451_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_2
XANTENNA__13469__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout541 _06382_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_4
Xfanout552 net553 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09705__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14130__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _06162_ _06163_ _06164_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__or4_1
Xfanout563 _04557_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout585 _04157_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12920_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] _07243_ net1031 vssd1 vssd1
+ vccd1 vccd1 _03618_ sky130_fd_sc_hd__mux2_1
Xfanout596 _03747_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12851_ net2479 net303 net368 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13661__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ net3042 net256 net480 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ net1174 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ net2475 net271 net375 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XANTENNA__11247__A3 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ net1407 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XANTENNA__08982__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11733_ net681 _07082_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11652__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12277__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17240_ clknet_leaf_28_wb_clk_i _02800_ _01103_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14452_ net1391 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
XANTENNA__16184__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14197__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11664_ net1934 net1158 net568 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1
+ vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08056__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _04903_ vssd1 vssd1
+ vccd1 vccd1 _03756_ sky130_fd_sc_hd__nand2_1
X_17171_ clknet_leaf_50_wb_clk_i _02731_ _01034_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10615_ _06414_ net523 vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__and2_1
X_14383_ net1329 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ net496 _07812_ net2755 net838 vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16122_ net1383 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ net23 net799 net594 net2990 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10546_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] net656 net629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__a22o_1
Xwire964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ net1355 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__inv_2
X_13265_ net93 net816 net600 net1953 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
X_10477_ _06738_ _06739_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__or3_1
XANTENNA__08503__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ net1279 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XANTENNA__12904__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ net2897 net279 net440 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
XANTENNA__09376__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ net2820 net2699 net819 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11183__A2 _07139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12147_ net2223 net219 net448 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12740__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14121__A2 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16955_ clknet_leaf_36_wb_clk_i _02515_ _00818_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12078_ net2746 net222 net457 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
X_15906_ net1345 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__inv_2
X_11029_ net538 _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__or2_1
XANTENNA__10143__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16886_ clknet_leaf_33_wb_clk_i _02446_ _00749_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15837_ net1281 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__inv_2
XANTENNA__10694__A1 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09053__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10199__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15768_ net1254 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__inv_2
XANTENNA__09988__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16527__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14719_ net1321 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
X_17507_ clknet_leaf_133_wb_clk_i _03067_ _01370_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12187__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15699_ net1187 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08240_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[116\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ net1038 vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
XANTENNA__14188__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17438_ clknet_leaf_3_wb_clk_i _02998_ _01301_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18116__1490 vssd1 vssd1 vccd1 vccd1 _18116__1490/HI net1490 sky130_fd_sc_hd__conb_1
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08171_ _04571_ _04572_ _04570_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a21oi_1
X_17369_ clknet_leaf_17_wb_clk_i _02929_ _01232_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11946__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17922__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_84_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_41_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09228__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_11_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08575__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12650__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__A3 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14112__A2 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17302__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ net579 _05888_ _05854_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout646_A _04751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1388_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _05815_ _05817_ _05819_ _05789_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a31o_2
XANTENNA__13623__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17452__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09260__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ net1079 net857 vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__and2_2
XFILLER_0_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12097__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _05747_ _05749_ _05750_ _05721_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_8_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14179__A2 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[31\] net752 net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12825__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08369_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] vssd1 vssd1 vccd1
+ vccd1 _04633_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _06662_ _06663_ net578 vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ _06777_ net332 vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ _06455_ _06594_ _06453_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13050_ net2400 net834 net354 _03686_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] _04487_ net766 _04719_ net1116
+ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09138__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11165__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13656__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ net495 _07845_ _08012_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10193_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] net962 vssd1
+ vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__and3_1
XANTENNA__12560__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10373__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1303 net1306 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__buf_4
XFILLER_0_44_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1314 net1338 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__buf_4
Xfanout1325 net1338 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__buf_2
XANTENNA__14103__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09435__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1336 net1337 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__buf_4
Xfanout1347 net1348 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__buf_4
Xfanout360 _03665_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_6
Xfanout1358 net1359 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__buf_4
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1369 net1370 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__buf_4
Xfanout371 _03571_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_6
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16740_ clknet_leaf_128_wb_clk_i _02300_ _00603_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout382 _03569_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_8
X_13952_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] net3226 vssd1 vssd1 vccd1
+ vccd1 _04145_ sky130_fd_sc_hd__nand2_1
Xfanout393 _03566_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
XFILLER_0_89_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08869__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13862__A1 team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ net366 _03604_ _03605_ net1056 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a32o_1
XANTENNA__11873__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16671_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[25\]
+ _00534_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13883_ _04505_ net1679 _03575_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_134_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11904__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15622_ net1275 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
X_12834_ net2656 net236 net367 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15553_ net1292 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
XANTENNA__09601__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12765_ net3164 net208 net377 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14504_ net1345 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17945__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11716_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _07856_ vssd1 vssd1
+ vccd1 vccd1 _07857_ sky130_fd_sc_hd__and2_1
X_15484_ net1234 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
X_12696_ _08008_ _08017_ net488 vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__and3_4
XFILLER_0_51_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17223_ clknet_leaf_126_wb_clk_i _02783_ _01086_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14435_ net1279 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12735__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09046__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11647_ team_01_WB.instance_to_wrap.cpu.DM0.enable net679 vssd1 vssd1 vccd1 vccd1
+ _07835_ sky130_fd_sc_hd__or2_2
XFILLER_0_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13420__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17154_ clknet_leaf_144_wb_clk_i _02714_ _01017_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
Xinput35 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XFILLER_0_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14366_ net1326 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
Xinput46 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
X_11578_ _04482_ _07794_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput57 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16105_ net1364 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__inv_2
Xhold808 team_01_WB.instance_to_wrap.cpu.c0.count\[12\] vssd1 vssd1 vccd1 vccd1 net2424
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13317_ net2905 net813 net807 net2135 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a22o_1
Xhold819 _04136_ vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] net721 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__a22o_1
X_17085_ clknet_leaf_130_wb_clk_i _02645_ _00948_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14297_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\] _04195_ net1912 vssd1
+ vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ net1410 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__inv_2
X_13248_ net52 net51 net54 net53 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09048__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15347__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13550__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17325__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__B1 _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ net3121 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\] net824 vssd1 vssd1
+ vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1508 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3124 sky130_fd_sc_hd__dlygate4sd3_1
X_17987_ clknet_leaf_57_wb_clk_i _03536_ _01807_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1519 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3135 sky130_fd_sc_hd__dlygate4sd3_1
X_16938_ clknet_leaf_43_wb_clk_i _02498_ _00801_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09521__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16869_ clknet_leaf_133_wb_clk_i _02429_ _00732_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11814__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] net618 _05663_
+ _05668_ _05669_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09341_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] net892 vssd1
+ vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09285__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08408__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15810__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__A1 _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09272_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[15\] net842 vssd1
+ vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_115_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _04502_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12645__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout227_A _07911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ net1736 net551 net348 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1
+ vccd1 vccd1 _03541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08424__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08796__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] team_01_WB.instance_to_wrap.cpu.f0.num\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1136_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08548__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_A _03747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12380__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1303_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09255__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08987_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] net867
+ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A2 _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__B _06992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout930_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09608_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] net896 vssd1
+ vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ net540 _06953_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] net850 vssd1
+ vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13072__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ net2703 net246 net403 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16992__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11501_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] _07741_ _07747_ vssd1 vssd1 vccd1
+ vccd1 _03373_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12481_ net2072 net278 net412 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XANTENNA__12555__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14336__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\] _04239_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\]
+ _04376_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__a221o_1
X_11432_ _04593_ _07683_ _07690_ net1162 vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__a22o_1
XANTENNA__09579__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10583__B team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08787__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16222__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\] _04263_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11363_ _04959_ _06935_ _06941_ net322 vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17348__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13102_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\] _06244_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10314_ _06575_ _06576_ _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__or3_1
XFILLER_0_132_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14082_ net789 _04232_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and3_4
X_11294_ _07465_ _07470_ net539 vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__mux2_1
X_13033_ _04954_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__o21a_1
X_17910_ clknet_leaf_101_wb_clk_i _03460_ _01730_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\]
+ sky130_fd_sc_hd__dfstp_1
X_10245_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\] net651 net646 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__a22o_1
XANTENNA__12290__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1100 net1105 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_1
XANTENNA__17498__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09165__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16372__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1111 net1113 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_2
X_10176_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\] net633 _06418_ _06422_
+ _06427_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09751__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__A1 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17841_ clknet_leaf_104_wb_clk_i _03391_ _01661_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_4
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_2
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_2
Xfanout1155 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1
+ net1155 sky130_fd_sc_hd__buf_2
Xfanout1166 net1167 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10104__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1177 net1179 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_4
X_17772_ clknet_leaf_95_wb_clk_i _03330_ _01593_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14984_ net1181 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
Xfanout190 _07874_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
Xfanout1188 net1194 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1199 net1203 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_4
X_16723_ clknet_leaf_22_wb_clk_i _02283_ _00586_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13935_ net1164 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[16\] sky130_fd_sc_hd__and3b_1
XFILLER_0_117_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13415__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16654_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[8\]
+ _00517_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13866_ team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] _04139_ _04140_ net1161 vssd1
+ vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08509__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15605_ net1176 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12817_ net2304 net265 net372 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
XANTENNA__09331__C net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16585_ clknet_leaf_86_wb_clk_i _02213_ _00448_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13797_ _07705_ _07784_ net484 vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15536_ net1264 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
XANTENNA__11074__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12748_ net2998 net246 net379 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15467_ net1206 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
X_12679_ net3112 net278 net388 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ clknet_leaf_32_wb_clk_i _02766_ _01069_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14418_ net1392 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18186_ net1560 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15398_ net1274 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08778__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17137_ clknet_leaf_24_wb_clk_i _02697_ _01000_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14349_ net2021 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold605 _03324_ vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold616 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net2232
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ clknet_leaf_48_wb_clk_i _02628_ _00931_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16019_ net1386 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__inv_2
XANTENNA__13523__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08910_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\] net873
+ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__and3_1
X_09890_ net1100 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\] net894 vssd1
+ vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12877__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10888__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\] net905
+ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09506__C net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1305 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net2932
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16865__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] net695 _05023_
+ _05027_ _05028_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__a2111o_1
Xhold1338 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1 vccd1
+ net2965 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11398__A_N _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13325__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08419__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1086_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09324_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\] net903
+ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12883__B _07640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09255_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\] net863 vssd1
+ vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout511_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12375__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1253_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout609_A _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _04568_ _04601_ _04602_ net553 net1659 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18139__1513 vssd1 vssd1 vccd1 vccd1 _18139__1513/HI net1513 sky130_fd_sc_hd__conb_1
XFILLER_0_105_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09186_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] net666 vssd1 vssd1
+ vccd1 vccd1 _05450_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08137_ team_01_WB.instance_to_wrap.cpu.K0.code\[2\] _04563_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__or3b_2
XFILLER_0_82_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10040__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_83_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08068_ team_01_WB.instance_to_wrap.cpu.f0.num\[3\] vssd1 vssd1 vccd1 vccd1 _04499_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout880_A _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17640__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10030_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[4\] net853 vssd1
+ vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17790__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ net2902 net220 net467 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13293__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13720_ _07681_ _04037_ _04039_ net783 net1627 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__o32a_1
X_10932_ net344 _07156_ _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10500__B1 _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17020__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13651_ _07495_ _03981_ net769 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10863_ _06778_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10297__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12602_ net2651 net203 net396 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
XANTENNA__15450__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16370_ clknet_leaf_104_wb_clk_i _02004_ _00238_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
X_13582_ net966 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _03922_ _03923_
+ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10794_ net549 _04828_ net500 vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08990__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15321_ net1190 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
X_12533_ net3208 net191 net403 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12285__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17170__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18040_ net1430 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_15252_ net1241 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
X_12464_ net2756 net213 net418 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16738__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14203_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\] _04249_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\]
+ _04358_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _06526_ vssd1 vssd1 vccd1
+ vccd1 _07678_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183_ net1248 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
X_12395_ net2597 net308 net426 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08999__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14134_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[9\] _04267_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[25\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11346_ _07001_ _07352_ _07609_ _07079_ _07608_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__a221o_1
XANTENNA__09972__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14065_ net792 net791 _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__and3_4
X_11277_ _05688_ net337 _06985_ _05686_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__o22a_1
XANTENNA__08511__B net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ net2908 net294 net362 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
X_10228_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] net843 vssd1
+ vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__and3_1
XANTENNA__09724__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09326__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_135_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08932__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17824_ clknet_leaf_80_wb_clk_i _03381_ _01645_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10159_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] net899 vssd1
+ vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__and3_1
Xhold2 team_01_WB.instance_to_wrap.a1.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 net1618
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11872__B _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17755_ clknet_leaf_115_wb_clk_i _03313_ _01576_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_14967_ net1243 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13284__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16706_ clknet_leaf_142_wb_clk_i _02266_ _00569_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11295__A1 _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13918_ net3268 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[31\]
+ sky130_fd_sc_hd__and2_1
X_17686_ clknet_leaf_75_wb_clk_i _03246_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14898_ net1188 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
XANTENNA__08160__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13849_ team_01_WB.instance_to_wrap.cpu.c0.count\[4\] _04111_ team_01_WB.instance_to_wrap.cpu.c0.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a21o_1
XANTENNA__09061__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16637_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[23\]
+ _00500_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14233__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17513__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09996__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16568_ clknet_leaf_13_wb_clk_i _02196_ _00431_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12195__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15519_ net1294 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16499_ clknet_leaf_101_wb_clk_i net2948 _00362_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09040_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\] net700 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10270__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18238_ net603 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17663__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18169_ net1543 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
Xhold402 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10558__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold413 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold424 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold435 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _03447_ vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08702__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[24\] vssd1 vssd1 vccd1 vccd1
+ net2084 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[5\] net916 vssd1
+ vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold479 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout904 net906 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08421__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09176__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout915 _04682_ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_6
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09715__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout926 _04668_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_8
X_09873_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\] _04641_ _04676_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__a22o_1
Xfanout937 net939 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_4
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_4
Xfanout959 net960 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__buf_4
Xhold1102 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\] vssd1 vssd1 vccd1 vccd1
+ net2718 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] net725 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a22o_1
Xhold1113 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 _03478_ vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09533__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11782__B _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1157 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\] net948 vssd1
+ vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout461_A _08015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] net616 net615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08151__B2 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12894__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout726_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1370_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15270__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09307_ _05568_ _05569_ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11303__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09238_ _05490_ _05499_ _05500_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11022__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] net748 net720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a22o_1
XANTENNA__12833__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10549__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ _06885_ net324 _07457_ _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__o31a_1
XFILLER_0_121_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net3205 net220 net444 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11131_ _06179_ _06601_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold980 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold991 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[94\] vssd1 vssd1 vccd1 vccd1
+ net2607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14160__B1 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13934__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _06033_ _06604_ _05760_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10013_ _06275_ _06276_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] net761
+ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__15445__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ net1396 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08985__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1350 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13266__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16410__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14752_ net1223 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17540_ clknet_leaf_139_wb_clk_i _03100_ _01403_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11964_ net2429 net293 net474 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13703_ _04466_ _04467_ _07719_ _04465_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17471_ clknet_leaf_2_wb_clk_i _03031_ _01334_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ _07177_ _07178_ net528 vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__mux2_1
X_14683_ net1363 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11895_ net678 _07121_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__nand2_1
XANTENNA_output109_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16422_ clknet_leaf_83_wb_clk_i _02050_ _00285_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13634_ _07344_ _03967_ net770 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__mux2_1
X_10846_ net511 _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17686__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16353_ clknet_leaf_73_wb_clk_i net1638 _00221_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13565_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _03909_ net1066 vssd1
+ vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
X_10777_ _07038_ _07040_ net512 vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__mux2_1
XANTENNA__08506__B net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15304_ net1181 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12516_ net2943 net277 net409 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ clknet_leaf_86_wb_clk_i _01918_ _00152_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13496_ _03847_ _03848_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15235_ net1225 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
X_18023_ net1417 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_23_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ net1931 net252 net417 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__mux2_1
XANTENNA__12743__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10004__A2 _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15166_ net1297 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12378_ net3104 net283 net425 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
X_14117_ net788 _04232_ _04241_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__and3_4
X_11329_ net525 _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__nand2_1
X_15097_ net1193 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
XANTENNA__17066__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14151__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ _04215_ net566 _04214_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09056__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12701__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11883__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17807_ clknet_leaf_68_wb_clk_i _03364_ _01628_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_18138__1512 vssd1 vssd1 vccd1 vccd1 _18138__1512/HI net1512 sky130_fd_sc_hd__conb_1
XFILLER_0_94_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15999_ net1388 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11094__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\] net943 vssd1
+ vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__and3_1
X_17738_ clknet_leaf_95_wb_clk_i _03296_ _01559_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\] net665 net663 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17669_ clknet_leaf_129_wb_clk_i _03229_ _01532_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08684__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10491__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__A0 _07033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08416__B net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09023_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\] net962 vssd1
+ vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and3_1
XANTENNA__13717__B1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12653__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1049_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[5\] vssd1 vssd1 vccd1 vccd1
+ net1826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09528__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 net84 vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 _01977_ vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold243 net113 vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _03298_ vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold265 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 net159 vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1216_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 _02072_ vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 net703 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_6
Xhold298 _01996_ vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 net714 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
XFILLER_0_1_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09925_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] net690 _06186_ _06187_
+ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__a2111o_1
Xfanout723 net724 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_6
Xfanout734 _04660_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
Xfanout745 _04648_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_6
XANTENNA_fanout676_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17559__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[6\] net927 vssd1
+ vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__and3_1
Xfanout767 _04626_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_2
Xfanout778 net780 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
Xfanout789 _04230_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09263__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\] net927 vssd1
+ vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09787_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\] net747 net730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout843_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08738_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] net631 _05001_
+ net670 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a211o_1
XANTENNA__10202__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _04921_ _04926_ _04930_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14609__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10700_ _06960_ _06963_ net525 vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11680_ net2033 net1160 net569 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _06600_ _06893_ _06892_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09624__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ net6 net799 net593 net3093 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] net666 _06816_ _06825_
+ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o22a_4
XFILLER_0_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13708__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12301_ net1975 net192 net427 vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
XANTENNA__11163__A1_N _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ net1839 net813 net599 team_01_WB.instance_to_wrap.a1.ADR_I\[10\] vssd1 vssd1
+ vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
XANTENNA__14344__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\] net661 net619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\]
+ _06756_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15020_ net1263 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
X_12232_ net2876 net211 net442 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_1
XANTENNA__09438__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09927__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12163_ net2872 net307 net450 vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A0 _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14133__B1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ _07375_ _07377_ _07374_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16971_ clknet_leaf_47_wb_clk_i _02531_ _00834_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12094_ net2057 net259 net457 vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11907__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11045_ _06832_ _06933_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__nand2_1
X_15922_ net1352 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16926__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ net1217 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__inv_2
XANTENNA__09604__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ net1362 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12996_ net2751 net226 net360 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
X_15784_ net1204 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__inv_2
XANTENNA__08115__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09312__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17523_ clknet_leaf_21_wb_clk_i _03083_ _01386_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11947_ net2395 net254 net472 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__mux2_1
X_14735_ net1314 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XANTENNA__12738__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14519__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13423__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14666_ net1409 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
X_17454_ clknet_leaf_52_wb_clk_i _03014_ _01317_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _07991_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__inv_2
XANTENNA__11670__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16405_ clknet_leaf_75_wb_clk_i _02033_ _00268_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_13617_ _03953_ _03952_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] net969
+ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a2bb2o_1
X_10829_ _06752_ _06807_ net498 vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17385_ clknet_leaf_38_wb_clk_i _02945_ _01248_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14597_ net1375 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16336_ clknet_leaf_62_wb_clk_i net1752 _00204_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
X_13548_ net185 _03893_ _03894_ net771 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a211o_1
XANTENNA__16306__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16267_ clknet_leaf_69_wb_clk_i _01904_ _00135_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12473__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13479_ _03830_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ clknet_leaf_83_wb_clk_i _03555_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_15218_ net1188 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XANTENNA__09918__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16198_ clknet_leaf_94_wb_clk_i _01865_ _00066_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12922__B2 _03619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ net1216 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
XANTENNA__16456__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09710_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] net928
+ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09083__A _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\] net926
+ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17851__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[8\] net745 net731 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08523_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\] net634 net623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\]
+ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a221o_1
XANTENNA__09811__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12648__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11110__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10464__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ _04629_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__or4_1
XANTENNA__11661__B2 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\] net963 vssd1
+ vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout424_A _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1166_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10216__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11413__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17231__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12383__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1333_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09006_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] net651 _05258_
+ _05259_ _05262_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09258__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14115__B1 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16949__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net524 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_2
XANTENNA__11727__S net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 net533 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_2
Xfanout542 net544 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
X_09908_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\] net658 _04777_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__a22o_1
Xfanout553 _04562_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 _04557_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_2
Xfanout586 net588 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_4
Xfanout597 net598 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_4
X_09839_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[7\] net608 _06075_ _06085_
+ _06090_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08896__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ net3034 net262 net368 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net775 _07926_ _07928_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12781_ net2460 net246 net376 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XANTENNA__12558__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14339__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18209__1583 vssd1 vssd1 vccd1 vccd1 _18209__1583/HI net1583 sky130_fd_sc_hd__conb_1
XANTENNA__13243__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14520_ net1411 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11732_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\] net674 net774 vssd1 vssd1
+ vccd1 vccd1 _07872_ sky130_fd_sc_hd__o21a_1
XANTENNA__11652__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14451_ net1391 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11663_ net1648 net1158 net567 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1
+ vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] _04903_ vssd1 vssd1
+ vccd1 vccd1 _03755_ sky130_fd_sc_hd__or2_1
XANTENNA__10207__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17170_ clknet_leaf_31_wb_clk_i _02730_ _01033_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10614_ _05281_ _05348_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__and2_1
X_14382_ net1328 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09073__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[29\] net572 vssd1 vssd1 vccd1
+ vccd1 _07812_ sky130_fd_sc_hd__nand2_1
X_16121_ net1387 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13333_ net25 net801 net596 net3218 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[24\] net644 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\]
+ _06808_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__a221o_1
XANTENNA__12293__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18137__1511 vssd1 vssd1 vccd1 vccd1 _18137__1511/HI net1511 sky130_fd_sc_hd__conb_1
XFILLER_0_24_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16052_ net1410 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13264_ net1786 net816 net600 team_01_WB.instance_to_wrap.a1.ADR_I\[27\] vssd1 vssd1
+ vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
X_10476_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\] net734 net717 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15003_ net1298 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_12215_ net2042 net251 net441 vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13195_ net1732 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] net824 vssd1 vssd1
+ vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12146_ net2887 net282 net449 vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17874__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16954_ clknet_leaf_36_wb_clk_i _02514_ _00817_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12077_ net2773 net226 net455 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15905_ net1349 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__inv_2
X_11028_ _07131_ _07232_ net520 vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__mux2_1
XANTENNA__09334__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16885_ clknet_leaf_25_wb_clk_i _02445_ _00748_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08887__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17104__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15836_ net1270 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09631__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12979_ net365 _03659_ _03660_ net1053 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15767_ net1239 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
XANTENNA__12468__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17506_ clknet_leaf_143_wb_clk_i _03066_ _01369_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14718_ net1411 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XANTENNA__10446__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15698_ net1184 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17437_ clknet_leaf_127_wb_clk_i _02997_ _01300_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14649_ net1402 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_16 net2932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08170_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[5\] team_01_WB.instance_to_wrap.cpu.K0.code\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__or4b_2
XANTENNA__13396__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17368_ clknet_leaf_28_wb_clk_i _02928_ _01231_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16319_ clknet_leaf_74_wb_clk_i _01953_ _00187_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17299_ clknet_leaf_50_wb_clk_i _02859_ _01162_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_113_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__15808__A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__14712__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__09525__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09524__B1 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout374_A _03571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09624_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] net669 _05882_ _05887_
+ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_39_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09541__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _05808_ _05809_ _05810_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__nor4_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12378__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A _06382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08506_ net1001 net846 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__and2_2
XANTENNA__10437__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _05739_ _05740_ _05741_ _05742_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__or4_2
XFILLER_0_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08437_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[31\] net732 net698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\]
+ _04654_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout806_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17747__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13387__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ net1155 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 _04632_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ net3188 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\] net1049 vssd1 vssd1
+ vccd1 vccd1 _03448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10070__B1 _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13002__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10330_ _06525_ _06593_ _06524_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17897__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12841__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _06485_ net517 vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12898__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ net3185 net210 net468 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ _06453_ _06454_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__or2_1
XANTENNA__10373__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 net1306 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__buf_2
Xfanout1315 net1316 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__buf_4
Xfanout1326 net1327 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__buf_4
Xfanout1337 net1338 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout350 _03751_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xfanout1348 net1349 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__clkbuf_4
Xfanout361 _03665_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_4
XANTENNA__09515__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1359 net1360 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__clkbuf_4
Xfanout372 _03571_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_4
X_13951_ net1617 net1169 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.next_keyvalid
+ sky130_fd_sc_hd__nor2_1
Xfanout383 _03568_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_8
Xfanout394 _03566_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08869__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15453__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] vssd1 vssd1 vccd1
+ vccd1 _03605_ sky130_fd_sc_hd__or2_2
XFILLER_0_57_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16670_ clknet_leaf_113_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[24\]
+ _00533_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13882_ _04505_ net3090 team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] _07834_ vssd1
+ vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__a22o_1
XANTENNA__17277__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15621_ net1233 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
X_12833_ net1999 net203 net367 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XANTENNA__13075__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12288__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10428__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ net3157 net190 net375 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15552_ net1252 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14503_ net1343 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
X_11715_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\]
+ _07855_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15483_ net1299 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ net2497 net213 net390 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11920__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13701__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17222_ clknet_leaf_139_wb_clk_i _02782_ _01085_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14434_ net1234 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XANTENNA__13378__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11646_ team_01_WB.instance_to_wrap.cpu.DM0.enable net679 vssd1 vssd1 vccd1 vccd1
+ _07834_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1326 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XANTENNA__13420__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17153_ clknet_leaf_137_wb_clk_i _02713_ _01016_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_1
Xinput36 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
XFILLER_0_128_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _07800_ _07798_ vssd1 vssd1 vccd1
+ vccd1 _03350_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput47 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13316_ net1698 net811 net805 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\] vssd1
+ vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a22o_1
Xinput58 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_16104_ net1377 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__inv_2
Xinput69 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10528_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[24\] net956
+ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__and3_1
X_17084_ clknet_leaf_15_wb_clk_i _02644_ _00947_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold809 team_01_WB.instance_to_wrap.cpu.f0.num\[30\] vssd1 vssd1 vccd1 vccd1 net2425
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ net1980 _04195_ _04442_ net1367 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09329__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13247_ _03728_ _03729_ _03730_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16035_ net1401 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12751__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12889__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ _06668_ _06721_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13550__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09626__A _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13178_ net2075 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\] net818 vssd1 vssd1
+ vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
X_18240__1593 vssd1 vssd1 vccd1 vccd1 _18240__1593/HI net1593 sky130_fd_sc_hd__conb_1
X_12129_ net2503 net311 net454 vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17986_ clknet_leaf_64_wb_clk_i _03535_ _01806_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1509 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3125 sky130_fd_sc_hd__dlygate4sd3_1
X_16937_ clknet_leaf_40_wb_clk_i _02497_ _00800_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09064__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16868_ clknet_leaf_128_wb_clk_i _02428_ _00731_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09361__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15819_ net1205 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__inv_2
XANTENNA__12198__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ clknet_leaf_0_wb_clk_i _02359_ _00662_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_09340_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] net863
+ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10419__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09285__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\] net856 vssd1
+ vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _04615_ _04616_ _04606_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13369__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08705__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08153_ net1882 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1
+ vccd1 vccd1 _03542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08424__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] _04494_ team_01_WB.instance_to_wrap.cpu.f0.num\[6\]
+ _04479_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12661__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1031_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1129_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09536__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18208__1582 vssd1 vssd1 vccd1 vccd1 _18208__1582/HI net1582 sky130_fd_sc_hd__conb_1
XFILLER_0_41_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout491_A _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A _03585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net1003 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\] net864
+ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__and3_1
XANTENNA__16174__CLK clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18136__1510 vssd1 vssd1 vccd1 vccd1 _18136__1510/HI net1510 sky130_fd_sc_hd__conb_1
XFILLER_0_93_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\] net881 vssd1
+ vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09702__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09538_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] net907 vssd1
+ vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__and3_1
XANTENNA__09276__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09469_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[12\] net868 vssd1
+ vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__and3_1
XANTENNA__12836__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11500_ team_01_WB.instance_to_wrap.cpu.f0.i\[25\] _07743_ vssd1 vssd1 vccd1 vccd1
+ _07747_ sky130_fd_sc_hd__nand2_1
XANTENNA__13521__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12480_ net2487 net250 net413 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] _07689_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13780__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14150_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\] _04227_ _04238_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\]
+ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__a22o_1
XANTENNA__14309__B1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ _04959_ _06838_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ net1701 net837 net357 _03720_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[0\] net748 _04672_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__and2b_2
XANTENNA__12571__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10880__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ _05962_ net343 _06988_ _05961_ _07556_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13032_ net2288 net834 net354 _03674_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08988__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[1\] net660 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a22o_1
XANTENNA_input52_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1103 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
X_17840_ clknet_leaf_88_wb_clk_i team_01_WB.instance_to_wrap.cpu.f0.next_write_i _01660_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_i sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10175_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[2\] net866 vssd1
+ vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__and3_1
XANTENNA__10897__A2 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1123 net1140 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_4
Xfanout1134 net1140 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1145 net1146 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_2
Xfanout1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\] vssd1 vssd1 vccd1 vccd1
+ net1156 sky130_fd_sc_hd__clkbuf_4
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_2
X_17771_ clknet_leaf_95_wb_clk_i _03329_ _01592_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14983_ net1180 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
Xfanout191 _07874_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16667__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1189 net1194 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_4
XANTENNA__11915__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16722_ clknet_leaf_23_wb_clk_i _02282_ _00585_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13934_ net1164 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[15\] sky130_fd_sc_hd__and3b_1
XANTENNA__11846__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17912__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16653_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[7\]
+ _00516_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09612__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ team_01_WB.instance_to_wrap.cpu.DM0.state\[1\] team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08509__B net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ net1241 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
X_12816_ net2012 net269 net373 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XANTENNA__10120__A _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16584_ clknet_leaf_72_wb_clk_i _02212_ _00447_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13796_ net1805 net782 _04096_ _04098_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14260__A2 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ net1269 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ net3115 net274 net382 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
XANTENNA__12746__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14527__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12678_ net2106 net250 net389 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
X_15466_ net1197 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17205_ clknet_leaf_26_wb_clk_i _02765_ _01068_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14417_ net1309 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
X_11629_ net1861 net839 _07808_ _07829_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__o22a_1
X_18185_ net1559 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15397_ net1225 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08778__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17136_ clknet_leaf_24_wb_clk_i _02696_ _00999_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13771__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14348_ net1716 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09059__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold606 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold617 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ clknet_leaf_46_wb_clk_i _02627_ _00930_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12481__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold639 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[26\] vssd1 vssd1 vccd1 vccd1
+ net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10790__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ net791 net790 net788 net1404 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__a31o_1
XANTENNA__13523__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ net1394 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire557_A _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17442__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11097__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\] net893 vssd1
+ vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1306 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1317 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net2933 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[22\] net749 _05017_
+ _05024_ _05026_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13287__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17969_ clknet_leaf_79_wb_clk_i team_01_WB.instance_to_wrap.cpu.f0.next_lcd_en _01789_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.enable sky130_fd_sc_hd__dfrtp_1
Xhold1328 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11825__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09091__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08419__B net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14251__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\] net881 vssd1
+ vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12656__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout337_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1079_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[15\] net860 vssd1
+ vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10684__B _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08205_ _04482_ _04566_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] net576 net577 vssd1 vssd1
+ vccd1 vccd1 _05449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1246_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ team_01_WB.instance_to_wrap.cpu.K0.code\[1\] team_01_WB.instance_to_wrap.cpu.K0.code\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08067_ team_01_WB.instance_to_wrap.cpu.f0.num\[4\] vssd1 vssd1 vccd1 vccd1 _04498_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12391__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1413_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout873_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17935__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13278__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[19\] net745 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11735__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ net1937 net282 net469 vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10931_ _06874_ _07159_ _07160_ _07192_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__o311a_1
XFILLER_0_98_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09432__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ _06832_ _06933_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__or2_1
X_13650_ _07968_ _03980_ net187 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12601_ net2739 net238 net395 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_13581_ net773 _07287_ net967 vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12566__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _04854_ net340 net339 _04852_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10875__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15320_ net1254 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
X_12532_ net2098 net194 net405 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ net2666 net290 net416 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
X_15251_ net1186 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _07677_ _07675_ vssd1
+ vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__mux2_1
X_14202_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\] _04255_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__a221o_1
X_15182_ net1230 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12394_ net2466 net313 net426 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14133_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\] _04233_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\]
+ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a22o_1
X_11345_ net545 _07364_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14064_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__and2_2
X_11276_ _05757_ _06905_ _06867_ _06856_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09607__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ net1898 net307 net363 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XANTENNA__09185__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10227_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] net903 vssd1
+ vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17823_ clknet_leaf_89_wb_clk_i _03380_ _01644_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10158_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] net852 vssd1
+ vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__and3_1
XANTENNA__13269__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 _02006_ vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13426__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17754_ clknet_leaf_114_wb_clk_i _03312_ _01575_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_10089_ net1103 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] net880 vssd1
+ vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14966_ net1303 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16705_ clknet_leaf_132_wb_clk_i _02265_ _00568_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13917_ net3271 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[30\]
+ sky130_fd_sc_hd__and2_1
X_17685_ clknet_leaf_74_wb_clk_i _03245_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09342__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11295__A2 _07555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14897_ net1246 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
X_16636_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[22\]
+ _00499_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13848_ net2459 _04121_ _04132_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[16\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14233__A2 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16567_ clknet_leaf_37_wb_clk_i _02195_ _00430_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12476__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18207__1581 vssd1 vssd1 vccd1 vccd1 _18207__1581/HI net1581 sky130_fd_sc_hd__conb_1
X_13779_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] net1065 _07707_ _04558_ vssd1
+ vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15518_ net1316 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16498_ clknet_leaf_102_wb_clk_i net2525 _00361_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17808__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ net603 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
X_15449_ net1190 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10007__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18168_ net1542 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11215__A_N _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09412__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\] vssd1 vssd1 vccd1 vccd1
+ net2019 sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ clknet_leaf_0_wb_clk_i _02679_ _00982_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold414 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold436 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ net1473 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17958__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold447 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09086__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold469 _02048_ vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[5\] net965 vssd1
+ vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__buf_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout927 _04666_ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_8
X_09872_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] net740 net728 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a22o_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_4
Xfanout949 _04650_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09814__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1103 _02102_ vssd1 vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ _05084_ _05085_ _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__or3_1
Xhold1114 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1125 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\] vssd1 vssd1 vccd1 vccd1
+ net2741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] net745 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a22o_1
Xhold1158 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09479__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08685_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\] net645 net622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a22o_1
XANTENNA__08687__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09252__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17338__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_A _08018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10494__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12894__B _07653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14224__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12386__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1363_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[14\] net724 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout719_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09651__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\] net741 net724 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[15\]
+ _05492_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13735__A1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[16\] net749 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout990_A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08119_ _04470_ team_01_WB.instance_to_wrap.cpu.f0.num\[18\] team_01_WB.instance_to_wrap.cpu.f0.num\[7\]
+ _04478_ _04547_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08611__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] net750 net719 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13010__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ net544 _07393_ _07392_ _07385_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09427__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold992 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[59\] vssd1 vssd1 vccd1 vccd1
+ net2608 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _05760_ _06033_ _06604_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10012_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ net1350 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ net1221 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XANTENNA__08678__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ net2591 net294 net474 vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09162__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13702_ net564 _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__nand2_1
XANTENNA__10485__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17470_ clknet_leaf_3_wb_clk_i _03030_ _01333_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ _07008_ _07013_ net512 vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__mux2_1
X_14682_ net1409 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
X_11894_ net2896 net290 net480 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux2_1
XANTENNA__14215__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16421_ clknet_leaf_75_wb_clk_i net3177 _00284_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10845_ _06347_ _06414_ net506 vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__mux2_1
X_13633_ _07954_ _03966_ net188 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__mux2_1
XANTENNA__12296__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16352_ clknet_leaf_66_wb_clk_i net1833 _00220_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08075__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ net767 _03907_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__a21boi_1
X_10776_ _07039_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15303_ net1182 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12515_ net1949 net216 net407 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16283_ clknet_leaf_85_wb_clk_i _01917_ _00151_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13495_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05167_ vssd1 vssd1
+ vccd1 vccd1 _03848_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18022_ net1416 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
X_12446_ net1888 net256 net416 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
X_15234_ net1290 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
XANTENNA__08803__A _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15165_ net1282 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ net3248 net224 net425 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14116_ net793 _04226_ _04243_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__and3_4
X_11328_ _06958_ _06974_ net514 vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__mux2_1
X_15096_ net1258 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
XANTENNA__09337__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14047_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] _04213_ vssd1 vssd1 vccd1
+ vccd1 _04215_ sky130_fd_sc_hd__and2_1
X_11259_ _05622_ _05756_ _07203_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18012__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16235__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17806_ clknet_leaf_59_wb_clk_i _03363_ _01627_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15998_ net1388 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17737_ clknet_leaf_96_wb_clk_i _03295_ _01558_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_14949_ net1232 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10476__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08470_ net1081 net903 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17668_ clknet_leaf_138_wb_clk_i _03228_ _01531_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14206__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16619_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[5\]
+ _00482_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17599_ clknet_leaf_5_wb_clk_i _03159_ _01462_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire889_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10779__A1 _07042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09022_ net1131 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] net957
+ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__and3_1
XANTENNA__17780__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09809__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold200 net129 vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold211 net87 vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10454__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout202_A _07888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 _02001_ vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08432__B net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 team_01_WB.instance_to_wrap.a1.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 net1849
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10400__A0 _06662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold244 _01965_ vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12940__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17010__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 team_01_WB.instance_to_wrap.cpu.f0.write_data\[21\] vssd1 vssd1 vccd1 vccd1
+ net1882 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16158__RESET_B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold277 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold288 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[126\] vssd1 vssd1 vccd1 vccd1
+ net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 net77 vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_4
X_09924_ net1136 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\] net939 vssd1
+ vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__and3_1
Xfanout713 net714 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_8
Xfanout724 _04669_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_8
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1111_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1209_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net737 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout746 _04646_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_8
X_09855_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] net938 vssd1
+ vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__and3_1
Xfanout757 net758 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_A _07804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _04626_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_2
Xfanout779 net780 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13066__A _05414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _05066_ _05067_ _05015_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or3b_1
X_09786_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] net918 vssd1
+ vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[23\] net664 net656 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08668_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[28\] net740 net716 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\]
+ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09872__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09710__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] net945
+ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13005__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ _06277_ net544 vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09624__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _06818_ _06820_ _06822_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12844__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net2117 net196 net429 vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XANTENNA__13708__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13280_ net1915 net812 net598 team_01_WB.instance_to_wrap.a1.ADR_I\[11\] vssd1 vssd1
+ vccd1 vccd1 _01994_ sky130_fd_sc_hd__a22o_1
X_10492_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[25\] net634 _04767_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _06756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231_ net3045 net292 net442 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09388__A1 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12162_ net3096 _07994_ net450 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10942__A1 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16258__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ net321 _07321_ _07376_ _07106_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16970_ clknet_leaf_42_wb_clk_i _02530_ _00833_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12093_ net1779 net298 net457 vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__mux2_1
X_18206__1580 vssd1 vssd1 vccd1 vccd1 _18206__1580/HI net1580 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08996__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ _05070_ _06613_ _06614_ _06833_ _05209_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__o2111ai_1
X_15921_ net1352 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15852_ net1264 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14803_ net1362 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XANTENNA__17653__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15783_ net1184 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
X_12995_ net2196 net200 net360 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11923__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17522_ clknet_leaf_31_wb_clk_i _03082_ _01385_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14734_ net1318 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11946_ net2323 net219 net472 vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09863__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13423__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17453_ clknet_leaf_19_wb_clk_i _03013_ _01316_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14665_ net1399 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _07848_ _07990_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ clknet_leaf_103_wb_clk_i _02032_ _00267_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13616_ net772 _07223_ net969 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a21o_1
X_17384_ clknet_leaf_62_wb_clk_i _02944_ _01247_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ _06643_ _06697_ net499 vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__mux2_1
XANTENNA__09615__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ net1399 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16335_ clknet_leaf_61_wb_clk_i _01969_ _00203_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_13547_ _07862_ _07894_ _07669_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o21a_1
XANTENNA__12754__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ _06843_ net346 _06871_ _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__a31o_2
XFILLER_0_54_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09629__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16266_ clknet_leaf_69_wb_clk_i _01903_ _00134_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17033__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08533__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13478_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _05380_ vssd1 vssd1
+ vccd1 vccd1 _03831_ sky130_fd_sc_hd__or2_1
X_18005_ clknet_leaf_82_wb_clk_i _03554_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_15217_ net1189 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
X_12429_ net1834 net294 net422 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
X_16197_ clknet_leaf_92_wb_clk_i _01864_ _00065_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12922__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13580__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ net1252 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
XANTENNA__09067__C net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10933__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15079_ net1180 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09364__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10697__A0 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\] net917 vssd1
+ vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__and3_1
XANTENNA__10303__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18095__1469 vssd1 vssd1 vccd1 vccd1 _18095__1469/HI net1469 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09571_ net1134 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] net928 vssd1
+ vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__and3_1
XANTENNA__11118__B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10449__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[31\] net657 net628 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a22o_1
XANTENNA__13614__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08453_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04629_ vssd1 vssd1 vccd1 vccd1
+ _04717_ sky130_fd_sc_hd__nor4_1
XFILLER_0_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09530__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08427__B net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08384_ net973 net961 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__and2_4
XFILLER_0_89_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11413__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12664__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1061_A team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09539__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__B _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09005_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[19\] net618 _05253_
+ _05254_ _05256_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16400__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1326_A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout510 _06523_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout521 net524 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_1
XANTENNA__09274__A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16550__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[6\] net649 _06170_ net673
+ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a211o_1
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_1
XANTENNA__17676__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09705__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout953_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _04202_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout576 _05243_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_4
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_2
X_09838_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\] net617 _06086_ _06092_
+ net672 vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__a2111o_1
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12839__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _05961_ _06032_ _06031_ _05892_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net681 _07243_ _07927_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12780_ net2090 net276 net376 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__A1 _06995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11731_ _07866_ _07870_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14450_ net1392 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17056__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11662_ net1996 net1158 net568 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1
+ vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13401_ _03752_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _05065_ _05043_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__nand2b_1
X_14381_ net1328 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
Xwire900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_2
X_11593_ net496 _07811_ net2056 net838 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12574__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire933 _04663_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_2
X_16120_ net1377 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__inv_2
X_10544_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[24\] net637 net618 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__a22o_1
X_13332_ net26 net798 net593 net2550 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16051_ net1401 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13263_ net95 net816 net600 net1773 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
X_10475_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[25\] net752 _06725_ _06730_
+ _06734_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_27_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15002_ net1259 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
X_12214_ net2885 net257 net440 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__mux2_1
XANTENNA__12904__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13194_ net2125 net1902 net818 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ net2714 net222 net449 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10822__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12076_ net2649 net200 net455 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
X_16953_ clknet_leaf_16_wb_clk_i _02513_ _00816_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ _05069_ _05210_ _07289_ _07290_ net344 vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__a311o_1
X_15904_ net1345 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__inv_2
XANTENNA__10123__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16884_ clknet_leaf_6_wb_clk_i _02444_ _00747_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10143__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15835_ net1298 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__inv_2
XANTENNA__09912__A _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13617__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12749__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15766_ net1258 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__inv_2
X_12978_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[2\] net1035 vssd1 vssd1 vccd1
+ vccd1 _03660_ sky130_fd_sc_hd__or2_1
XANTENNA__13947__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09836__A2 _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17505_ clknet_leaf_136_wb_clk_i _03065_ _01368_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14717_ net1404 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ net2967 net310 net478 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_1
XANTENNA__12840__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15697_ net1196 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17436_ clknet_leaf_15_wb_clk_i _02996_ _01299_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14648_ net1401 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_17 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ clknet_leaf_9_wb_clk_i _02927_ _01230_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12484__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14579_ net1344 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
XANTENNA__17549__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16318_ clknet_leaf_72_wb_clk_i _01952_ _00186_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09359__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17298_ clknet_leaf_31_wb_clk_i _02858_ _01161_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16249_ clknet_leaf_70_wb_clk_i _01886_ _00117_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_3_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__08575__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput179 net603 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10382__A2 _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13328__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09623_ _05883_ _05884_ _05885_ _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__or4_2
XANTENNA__09822__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12659__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout367_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[9\] net622 _05790_ _05794_
+ _05799_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17079__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11095__A0 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ net1111 net1115 net1107 net1109 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__and4bb_2
X_09485_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\] net624 _05748_ net670
+ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a211o_1
XANTENNA__09260__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A _06383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1276_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\] net754 net716 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\]
+ _04694_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12394__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08367_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] net1156 net765 vssd1 vssd1
+ vccd1 vccd1 _04631_ sky130_fd_sc_hd__and3b_1
XFILLER_0_68_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout701_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09269__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08298_ net2726 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16916__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11311__B _07555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _06485_ net512 vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12898__A1 _07324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08566__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _06453_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10373__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__buf_4
Xfanout1316 net1325 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__clkbuf_4
Xfanout1327 net1338 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09435__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 _06980_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
Xfanout1338 net1415 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__buf_4
Xfanout351 _03751_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1349 net1414 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__buf_2
Xfanout362 _03665_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11039__A _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13950_ net1163 net1057 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[31\] sky130_fd_sc_hd__and3b_1
Xfanout373 _03571_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_6
Xfanout384 _03568_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_4
Xfanout395 _03565_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_6
XANTENNA__09732__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ net1025 _07611_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12569__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] _03581_ _04143_ team_01_WB.instance_to_wrap.cpu.RU0.next_dhit
+ net796 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__a311o_1
X_15620_ net1226 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12832_ net2231 net239 net370 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14272__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15551_ net1295 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12763_ net2604 net195 net377 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XANTENNA__11625__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16446__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14502_ net1344 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
X_11714_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _07854_ vssd1 vssd1
+ vccd1 vccd1 _07855_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15482_ net1305 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
X_12694_ net2126 net292 net389 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17221_ clknet_leaf_131_wb_clk_i _02781_ _01084_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14433_ net1233 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ net1823 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] net841 vssd1 vssd1
+ vccd1 vccd1 _03316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11389__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17152_ clknet_leaf_0_wb_clk_i _02712_ _01015_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14364_ net1328 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _07700_ _07796_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__nor2_1
XANTENNA__08083__A _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09451__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
X_18094__1468 vssd1 vssd1 vccd1 vccd1 _18094__1468/HI net1468 sky130_fd_sc_hd__conb_1
Xinput48 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16103_ net1368 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__inv_2
XANTENNA__17841__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ net1761 net809 net804 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\] vssd1
+ vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a22o_1
Xinput59 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17083_ clknet_leaf_32_wb_clk_i _02643_ _00946_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10527_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[24\] net741 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__a22o_1
X_14295_ _04195_ _04199_ net1980 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a21oi_1
X_16034_ net1394 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__inv_2
X_13246_ net43 net42 net45 net44 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__or4_2
X_10458_ _06719_ _06720_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_21_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12889__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08811__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12889__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08557__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177_ net1657 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\] net828 vssd1 vssd1
+ vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
X_10389_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\] net634 net629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10364__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17991__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12128_ net2691 net260 net453 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__mux2_1
X_17985_ clknet_leaf_59_wb_clk_i _03534_ _01805_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16936_ clknet_leaf_46_wb_clk_i _02496_ _00799_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12059_ net2105 net244 net460 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
XANTENNA__09642__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17221__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__B _07441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ clknet_leaf_119_wb_clk_i _02427_ _00730_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15818_ net1201 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__inv_2
X_16798_ clknet_leaf_13_wb_clk_i _02358_ _00661_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14263__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15749_ net1226 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17371__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__A0 _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\] net904 vssd1
+ vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and3_1
XANTENNA__08692__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16939__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08221_ _04611_ _04612_ _04613_ _04614_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17419_ clknet_leaf_51_wb_clk_i _02979_ _01282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08152_ net1678 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1
+ vccd1 vccd1 _03543_ sky130_fd_sc_hd__a22o_1
XANTENNA__11412__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13330__C net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ _04505_ net1162 vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__nand2_1
XANTENNA__08796__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08548__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_124_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1024_A _04484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08985_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] net907
+ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__and3_1
XANTENNA__09255__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12389__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1393_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16469__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout749_A _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] net867 vssd1
+ vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__and3_1
XANTENNA__08720__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13057__A1 _05133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14254__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11068__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\] net883 vssd1
+ vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__and3_1
XANTENNA__11306__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09468_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[12\] net877 vssd1
+ vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08419_ net972 net913 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09399_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\] net868 vssd1
+ vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13013__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11430_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\]
+ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[0\] _07688_ vssd1 vssd1 vccd1 vccd1
+ _07689_ sky130_fd_sc_hd__or4_1
XFILLER_0_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ _05280_ _07624_ _07622_ _07614_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__o211a_2
XANTENNA__08787__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10312_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[0\] net750 _06563_ _06565_
+ _06568_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__a2111o_1
X_13100_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[6\] _06174_ net1035 vssd1
+ vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__mux2_2
XFILLER_0_85_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11791__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14080_ net793 net790 _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__and3_4
X_11292_ _05960_ net337 net336 _05959_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11054__A1_N net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10880__B _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13031_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\] _03673_ net1028 vssd1
+ vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__mux2_1
X_10243_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\] net882 vssd1
+ vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17244__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\] net887 vssd1
+ vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__and3_1
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09165__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[21\] vssd1 vssd1 vccd1 vccd1
+ net1113 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10897__A3 _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1124 net1126 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_2
XANTENNA__13683__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1135 net1140 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_4
Xfanout1146 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1
+ net1146 sky130_fd_sc_hd__buf_4
X_17770_ clknet_leaf_95_wb_clk_i net1862 _01591_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14982_ net1293 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
Xfanout1157 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1157
+ sky130_fd_sc_hd__buf_2
Xfanout1168 team_01_WB.instance_to_wrap.a1.BUSY_O vssd1 vssd1 vccd1 vccd1 net1168
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__10104__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1179 net1185 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16721_ clknet_leaf_21_wb_clk_i _02281_ _00584_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout192 _07874_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
XANTENNA__09462__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13933_ net1168 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[14\] sky130_fd_sc_hd__and3b_1
XANTENNA__11846__A2 _07510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17394__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08711__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16652_ clknet_leaf_88_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[6\]
+ _00515_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13048__A1 _05009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864_ net1156 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] team_01_WB.instance_to_wrap.cpu.DM0.enable
+ _04629_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or4_1
XANTENNA__08078__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14245__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ net1187 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__B _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ net2426 net273 net371 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16583_ clknet_leaf_66_wb_clk_i _02211_ _00446_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ net563 _07775_ _04097_ net786 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a31o_1
XANTENNA__10120__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11931__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15534_ net1231 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XANTENNA__13712__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ net2692 net218 net382 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15465_ net1210 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
X_12677_ net2172 net254 net388 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17204_ clknet_leaf_5_wb_clk_i _02764_ _01067_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14416_ net1309 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18184_ net1558 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
X_11628_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[12\] _07806_ vssd1 vssd1 vccd1
+ vccd1 _07829_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15396_ net1224 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ clknet_leaf_54_wb_clk_i _02695_ _00998_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08778__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14347_ net2877 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire560 _05164_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_1
X_11559_ _07701_ _07770_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__nor2_1
XANTENNA__18015__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17066_ clknet_leaf_48_wb_clk_i _02626_ _00929_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09637__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08541__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14278_ net1676 net584 _04432_ net1170 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10990__C1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16017_ net1363 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__inv_2
X_13229_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ net826 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1307 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 net2923
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16611__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1318 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] net752 net715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[22\]
+ _05018_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a221o_1
X_17968_ clknet_leaf_100_wb_clk_i net1714 _01788_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[127\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1329 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\] vssd1 vssd1 vccd1 vccd1
+ net2945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13606__B _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16919_ clknet_leaf_24_wb_clk_i _02479_ _00782_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_17899_ clknet_leaf_80_wb_clk_i net2727 _01719_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13039__A1 _06716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12002__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17887__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14718__A net1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[14\] net877
+ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ net997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] net871 vssd1
+ vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17117__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_A _07897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ _04579_ _04586_ _04588_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__or4_2
X_09184_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] net761 _05446_ _05447_
+ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a22o_2
XFILLER_0_69_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08135_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] _04504_ net564 _04560_ _04561_
+ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12672__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ team_01_WB.instance_to_wrap.cpu.f0.num\[9\] vssd1 vssd1 vccd1 vccd1 _04497_
+ sky130_fd_sc_hd__inv_2
XANTENNA__17267__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11525__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1406_A net1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15284__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[19\] net718 net701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11289__A0 _07010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ _05159_ _05160_ _05161_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18093__1467 vssd1 vssd1 vccd1 vccd1 _18093__1467/HI net1467 sky130_fd_sc_hd__conb_1
XANTENNA__13008__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ _07175_ _07193_ net542 vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14227__B1 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10500__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _06721_ _07124_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12847__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ net1981 net206 net396 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13580_ net186 _03920_ _03921_ net773 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09654__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10792_ _04851_ net336 net333 _04853_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__a22o_1
XANTENNA__12982__A1_N _07441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12531_ _07845_ _08012_ net489 vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__and3_4
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15250_ net1178 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
X_12462_ net2406 net295 net418 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13678__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14201_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\] _04261_ _04280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\]
+ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__a22o_1
X_11413_ net770 net187 _07674_ _07676_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15181_ net1213 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
XANTENNA__12582__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ net2662 _07989_ net425 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08999__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\] _04253_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[113\]
+ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a22o_1
XANTENNA__12961__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09457__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11344_ _06955_ _07011_ _07054_ _06964_ _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14063_ net791 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__inv_2
XANTENNA__16634__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ _05760_ _07199_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__a21o_1
X_13014_ net3234 net312 net363 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10226_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\] net895 vssd1
+ vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11926__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17822_ clknet_leaf_66_wb_clk_i _03379_ _01643_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_10157_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] net906 vssd1
+ vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08932__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13269__B2 team_01_WB.instance_to_wrap.a1.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 team_01_WB.instance_to_wrap.a1.ADR_I\[25\] vssd1 vssd1 vccd1 vccd1 net1620
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09192__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16784__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[3\] net899 vssd1
+ vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13426__B _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17753_ clknet_leaf_114_wb_clk_i _03311_ _01574_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_14965_ net1173 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ net3270 net795 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[29\]
+ sky130_fd_sc_hd__and2_1
X_16704_ clknet_leaf_140_wb_clk_i _02264_ _00567_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_17684_ clknet_leaf_74_wb_clk_i _03244_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10131__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14896_ net1307 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XANTENNA__14218__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16635_ clknet_leaf_106_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[21\]
+ _00498_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13847_ team_01_WB.instance_to_wrap.cpu.c0.count\[16\] _04121_ _04126_ vssd1 vssd1
+ vccd1 vccd1 _04132_ sky130_fd_sc_hd__nand3_1
XANTENNA__12757__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13442__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16566_ clknet_leaf_36_wb_clk_i _02194_ _00429_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13778_ _04473_ _07776_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15517_ net1282 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12729_ _07841_ _08017_ net488 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16497_ clknet_leaf_85_wb_clk_i _02125_ _00360_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18236_ net601 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16164__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15448_ net1255 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ net1541 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
XANTENNA__12492__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ net1187 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10558__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 _03465_ vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ clknet_leaf_13_wb_clk_i _02678_ _00981_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09367__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ net1472 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_44_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold426 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 team_01_WB.instance_to_wrap.a1.ADR_I\[11\] vssd1 vssd1 vccd1 vccd1 net2064
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08702__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold459 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[56\] vssd1 vssd1 vccd1 vccd1
+ net2075 sky130_fd_sc_hd__dlygate4sd3_1
X_17049_ clknet_leaf_18_wb_clk_i _02609_ _00912_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_09940_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] net949 vssd1
+ vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__and3_1
XANTENNA__10306__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11507__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09176__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout906 _04733_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_4
X_09871_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[6\] net744 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__a22o_1
Xfanout917 net919 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_4
Xfanout928 _04666_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
Xfanout939 _04659_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
XANTENNA__11836__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] net753 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1104 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\] vssd1 vssd1 vccd1 vccd1
+ net2731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[22\] net928 vssd1
+ vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__and3_1
XANTENNA__09533__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1148 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[114\] vssd1 vssd1 vccd1 vccd1
+ net2775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15832__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08684_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\] net640 net608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a221o_1
XANTENNA__14209__B1 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13680__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12667__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14448__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A _08019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1189_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16507__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[14\] net684 _05555_
+ _05562_ _05565_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11443__B1 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout614_A _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09236_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[15\] net746 net742 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13735__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15279__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09167_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\] net917
+ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__and3_1
XANTENNA__10915__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14183__A _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11746__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ _04469_ team_01_WB.instance_to_wrap.cpu.f0.num\[19\] _04495_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\]
+ _04523_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09098_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[17\] net723 _05351_ _05356_
+ _05358_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_128_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09708__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout983_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 _04480_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold960 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net346 _07122_ _07308_ _07310_ _07323_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__a311o_4
Xhold993 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14160__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _06265_ _06269_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08127__B1 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ net1307 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
X_11962_ net2785 net309 net474 vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__mux2_1
XANTENNA__13671__A1 _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ net1061 _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09740__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _07005_ _07009_ net513 vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__mux2_1
XANTENNA__12577__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ net1402 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
X_11893_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] _04622_ _08002_ _08003_
+ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__a22o_2
XANTENNA__11481__S team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16420_ clknet_leaf_103_wb_clk_i net2085 _00283_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13632_ _03946_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__or2_1
X_10844_ _06071_ _06141_ _06211_ _06277_ net504 net517 vssd1 vssd1 vccd1 vccd1 _07108_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17432__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16351_ clknet_leaf_66_wb_clk_i net1886 _00219_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13563_ net771 _07611_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10775_ net505 _06591_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15302_ net1281 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
X_12514_ net2327 net280 net409 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16282_ clknet_leaf_87_wb_clk_i _00013_ _00150_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13494_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _05167_ vssd1 vssd1
+ vccd1 vccd1 _03847_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18021_ net1598 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ net1290 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
XANTENNA__15189__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12445_ net2157 _07925_ net416 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
XANTENNA__10825__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15164_ net1270 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08091__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ net2612 net226 net423 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
X_14115_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\] _04275_ _04276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[40\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a221o_1
X_11327_ _06840_ net342 net339 _04907_ _07590_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10126__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15095_ net1238 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
X_14046_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\] _04213_ vssd1 vssd1 vccd1
+ vccd1 _04214_ sky130_fd_sc_hd__or2_1
XANTENNA__14151__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _07344_ _07368_ _07480_ _07521_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12162__A1 _07994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\] net731 net720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11189_ net539 _07134_ _07234_ _06991_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__a211o_1
X_17805_ clknet_leaf_59_wb_clk_i _03362_ _01626_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15997_ net1355 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__inv_2
XANTENNA__13111__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14948_ net1224 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
X_17736_ clknet_leaf_96_wb_clk_i _03294_ _01557_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11673__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879_ net1315 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XANTENNA__12487__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17667_ clknet_leaf_119_wb_clk_i _03227_ _01530_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16618_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[4\]
+ _00481_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17598_ clknet_leaf_3_wb_clk_i _03158_ _01461_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16549_ clknet_leaf_40_wb_clk_i _02177_ _00412_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13900__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17925__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] net937 vssd1
+ vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18219_ net1587 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12925__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092__1466 vssd1 vssd1 vccd1 vccd1 _18092__1466/HI net1466 sky130_fd_sc_hd__conb_1
Xhold201 _01980_ vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 _02003_ vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09528__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 net76 vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _01998_ vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\] vssd1 vssd1 vccd1 vccd1
+ net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 net111 vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10036__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold267 net149 vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_01_WB.instance_to_wrap.cpu.f0.i\[17\] vssd1 vssd1 vccd1 vccd1 net1894
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09923_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\] net954 vssd1
+ vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__and3_1
XANTENNA__09825__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold289 _02142_ vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 _04683_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_8
XFILLER_0_106_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout714 _04678_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13350__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout397_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09854_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] net946 vssd1
+ vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__and3_1
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_8
Xfanout758 _04637_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1104_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
X_08805_ _05043_ _05065_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13066__B _07803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09263__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[7\] net958 vssd1
+ vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08736_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\] net655 net652 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10202__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17455__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11664__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout731_A _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\] net736 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout829_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\] net925
+ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11416__B1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14906__A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10560_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\] net640 net635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\]
+ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10491_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\] net641 net627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12230_ net3039 net295 net442 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09438__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12860__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ net2721 net260 net449 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A2 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ _07091_ _07115_ net534 vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__mux2_1
XANTENNA__14133__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net3054 net243 net457 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__mux2_1
Xhold790 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13341__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _07301_ _07306_ _07304_ _07291_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__or4b_4
X_15920_ net1352 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__inv_2
X_15851_ net1209 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14802_ net1344 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XANTENNA__15472__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15782_ net1281 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__inv_2
X_12994_ net2419 net286 net360 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1490 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09470__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14733_ net1321 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XANTENNA__09312__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17521_ clknet_leaf_22_wb_clk_i _03081_ _01384_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11655__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11945_ net2236 net284 net471 vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08520__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17452_ clknet_leaf_45_wb_clk_i _03012_ _01315_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14664_ net1402 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XANTENNA__08086__A team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11876_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\]
+ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 _07990_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16403_ clknet_leaf_100_wb_clk_i _02031_ _00266_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13615_ net188 _07940_ _03951_ net770 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17383_ clknet_leaf_123_wb_clk_i _02943_ _01246_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10827_ _07087_ _07090_ net528 vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__mux2_1
X_14595_ net1371 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ clknet_leaf_65_wb_clk_i net1629 _00202_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13546_ _03857_ _03858_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__xor2_1
X_10758_ _07004_ _07021_ _06951_ _07003_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__a211o_1
XANTENNA__08814__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ clknet_leaf_70_wb_clk_i net1895 _00133_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13477_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] _05380_ vssd1 vssd1
+ vccd1 vccd1 _03830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10689_ _06868_ _06952_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12907__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18004_ clknet_leaf_82_wb_clk_i _03553_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_15216_ net1250 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12428_ net3152 net309 net421 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09379__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16196_ clknet_leaf_92_wb_clk_i _01863_ _00064_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08587__A0 _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15147_ net1209 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17328__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ net2701 net259 net492 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10394__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078_ net1275 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
XANTENNA__13332__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _04204_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__13883__A1 _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__A1 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09570_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] net947 vssd1
+ vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13635__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10022__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08521_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[31\] net619 net613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[31\]
+ _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a221o_1
X_17719_ clknet_leaf_111_wb_clk_i _03279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09811__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11110__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13106__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12010__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ _04628_ _04635_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08383_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] net958
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13630__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout312_A _07994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1054_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] net658 _05252_ _05257_
+ _05261_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13020__C1 _07803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09258__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12680__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1221_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1319_A net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__A2 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13323__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net513 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09906_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\] net641 net633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout522 net524 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout544 _06315_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
Xfanout566 _04202_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_1
Xfanout577 _05242_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
X_09837_ _06097_ _06098_ _06099_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or4_2
Xfanout588 _03585_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout599 _03742_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_4
XANTENNA_fanout946_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09768_ _05960_ _06029_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09290__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _04972_ _04980_ _04981_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _05923_ _05959_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13016__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11730_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _07865_ vssd1 vssd1
+ vccd1 vccd1 _07870_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11661_ net1782 net1158 net569 net1142 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12855__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _04850_ vssd1 vssd1
+ vccd1 vccd1 _03753_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ _05205_ _06873_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__o21ai_1
X_14380_ net1328 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[30\] net572 vssd1 vssd1 vccd1
+ vccd1 _07811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire912 _04728_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_144_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13331_ net1163 net801 team_01_WB.instance_to_wrap.a1.prev_BUSY_O vssd1 vssd1 vccd1
+ vccd1 _03748_ sky130_fd_sc_hd__or3b_1
XANTENNA__16225__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] net759 _06805_ _06806_
+ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__a22o_2
XFILLER_0_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16050_ net1405 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ net1808 net816 net600 team_01_WB.instance_to_wrap.a1.ADR_I\[29\] vssd1 vssd1
+ vccd1 vccd1 _02012_ sky130_fd_sc_hd__a22o_1
X_10474_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] net750 net747 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08569__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15001_ net1190 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12213_ net3229 net221 net439 vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12590__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\] net2101 net828 vssd1 vssd1
+ vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10376__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ net2592 net226 net447 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__mux2_1
XANTENNA__09465__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12117__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13314__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16952_ clknet_leaf_25_wb_clk_i _02512_ _00815_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12075_ net3123 net287 net455 vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11026_ _05210_ _07289_ _05069_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__a21oi_1
X_15903_ net1339 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__inv_2
XANTENNA__11876__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16883_ clknet_leaf_50_wb_clk_i _02443_ _00746_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08741__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ net1267 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08642__A_N _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13617__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18091__1465 vssd1 vssd1 vccd1 vccd1 _18091__1465/HI net1465 sky130_fd_sc_hd__conb_1
XANTENNA__09631__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ net1027 _07456_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nand2_1
X_15765_ net1177 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
X_17504_ clknet_leaf_141_wb_clk_i _03064_ _01367_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11235__A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14716_ net1408 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
X_11928_ net2423 net311 net477 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15696_ net1262 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17435_ clknet_leaf_37_wb_clk_i _02995_ _01298_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14647_ net1363 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _07849_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12765__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ clknet_leaf_30_wb_clk_i _02926_ _01229_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14578_ net1362 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XANTENNA__08544__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16317_ clknet_leaf_76_wb_clk_i _01951_ _00185_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
X_13529_ net771 _03878_ net1066 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__o21ai_1
X_17297_ clknet_leaf_21_wb_clk_i _02857_ _01160_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17150__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16248_ clknet_leaf_79_wb_clk_i _01885_ _00116_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16718__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XANTENNA_max_cap911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
X_16179_ clknet_leaf_90_wb_clk_i _01847_ _00047_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__10367__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10017__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12005__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16868__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08732__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[8\] net626 _05858_ _05864_
+ _05867_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13608__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09553_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] net639 _05816_ net671
+ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09541__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ net998 net877 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__and2_2
XANTENNA__11095__A1 _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09484_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] net660 net642 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[31\] net743 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a22o_1
XANTENNA__16248__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1269_A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\] _04629_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor3b_1
XANTENNA__08454__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08799__B1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ net2945 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] net1051 vssd1 vssd1
+ vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10070__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout896_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13544__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10190_ _06414_ net530 vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__nor2_1
XANTENNA__09763__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1306 net1307 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__buf_2
Xfanout1317 net1319 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__buf_4
XFILLER_0_100_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17793__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1328 net1329 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__buf_4
Xfanout330 _06990_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_4
Xfanout1339 net1349 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__buf_4
Xfanout341 _06980_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
Xfanout352 _03751_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09515__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11039__B _06867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 _03665_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_4
Xfanout374 _03571_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
Xfanout385 _03568_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
X_12900_ net2882 net607 net589 _03603_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a22o_1
XANTENNA__08723__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 _03565_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_4
X_13880_ net1165 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\] vssd1 vssd1 vccd1
+ vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_ihit sky130_fd_sc_hd__and2b_1
XFILLER_0_97_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12831_ net2698 net206 net370 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XANTENNA__13075__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ net1297 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XANTENNA__11086__A1 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12762_ _07842_ _08011_ net488 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__and3_4
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ net1344 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\]
+ _07853_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__and3_1
X_15481_ net1191 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12693_ net2557 net297 net390 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__mux2_1
XANTENNA__12585__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17173__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14432_ net1230 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
X_17220_ clknet_leaf_128_wb_clk_i _02780_ _01083_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11644_ net2741 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[1\] net841 vssd1 vssd1
+ vccd1 vccd1 _03317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17151_ clknet_leaf_1_wb_clk_i _02711_ _01014_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14363_ net1382 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
X_11575_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _07798_ _07799_ _07731_ vssd1 vssd1
+ vccd1 vccd1 _03351_ sky130_fd_sc_hd__a22o_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XFILLER_0_25_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16102_ net1371 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__inv_2
X_13314_ net109 net815 net806 net1700 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a22o_1
Xinput38 wb_rst_i vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_17082_ clknet_leaf_34_wb_clk_i _02642_ _00945_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput49 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_2
X_10526_ net971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\] net924 vssd1
+ vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14294_ _04195_ _04199_ _04441_ net1367 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_29_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11929__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16033_ net1365 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__inv_2
X_13245_ net70 net69 net41 net40 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10457_ _06719_ _06720_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09195__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09754__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ net2805 net2713 net826 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XANTENNA__08303__S net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] net665 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[27\]
+ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08962__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A2 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net2271 net298 net454 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10134__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17984_ clknet_leaf_61_wb_clk_i _03533_ _01804_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09923__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ net2599 net316 net461 vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
X_16935_ clknet_leaf_120_wb_clk_i _02495_ _00798_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08714__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net522 _06992_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__nor2_1
XANTENNA__13445__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16866_ clknet_leaf_144_wb_clk_i _02426_ _00729_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08539__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15817_ net1213 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
XANTENNA__09361__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16797_ clknet_leaf_130_wb_clk_i _02357_ _00660_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15748_ net1226 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10300__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10824__A1 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15679_ net1294 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08220_ _04607_ _04608_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__or4_2
X_17418_ clknet_leaf_43_wb_clk_i _02978_ _01281_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08151_ net1831 net551 net348 net1062 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09978__C1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11412__B _07441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08705__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17349_ clknet_leaf_133_wb_clk_i _02909_ _01212_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10309__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08082_ _04505_ net1162 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11001__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09536__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[19\] net861
+ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1017_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17046__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout477_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09605_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[8\] net850 vssd1
+ vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09271__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout644_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17196__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15570__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ net1015 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] net848 vssd1
+ vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09467_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\] net891 vssd1
+ vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout811_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14186__A _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08418_ net1147 net1154 net1151 net1150 vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] net885
+ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\] net1866 net1043 vssd1 vssd1
+ vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10043__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11360_ _06924_ net323 _07228_ _07623_ net345 vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__o32a_1
XFILLER_0_61_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08912__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10311_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] _04662_ net726 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ net535 _07462_ _07554_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18090__1464 vssd1 vssd1 vccd1 vccd1 _18090__1464/HI net1464 sky130_fd_sc_hd__conb_1
X_13030_ _04902_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o21a_1
X_10242_ net1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\] net907 vssd1
+ vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__and3_1
XANTENNA__14190__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13937__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13249__B net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\] net861 vssd1
+ vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__and3_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1114 net1116 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09743__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1136 net1140 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input38_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14981_ net1225 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
Xfanout1158 team_01_WB.instance_to_wrap.cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1158
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__16413__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16720_ clknet_leaf_24_wb_clk_i _02280_ _00583_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout193 _07874_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_1
X_13932_ net1167 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[13\] sky130_fd_sc_hd__and3b_1
XANTENNA__10503__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16651_ clknet_leaf_88_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[5\]
+ _00514_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13863_ _03744_ _04011_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15602_ net1178 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12814_ net2453 net246 net371 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16582_ clknet_leaf_66_wb_clk_i _02210_ _00445_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13794_ _04474_ _07774_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__C _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15533_ net1216 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
X_12745_ net2615 net279 net379 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ net1182 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
X_12676_ net2661 net219 net388 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12559__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17203_ clknet_leaf_21_wb_clk_i _02763_ _01066_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14415_ net1308 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11627_ net2810 net840 _07808_ _07828_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__o22a_1
X_18183_ net1557 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
X_15395_ net1223 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XANTENNA__10129__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17134_ clknet_leaf_51_wb_clk_i _02694_ _00997_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14346_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[12\] vssd1 vssd1 vccd1
+ vccd1 _02252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11231__A1 _06869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ team_01_WB.instance_to_wrap.cpu.f0.i\[8\] _07745_ _07786_ vssd1 vssd1 vccd1
+ vccd1 _03356_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09975__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire561 _05062_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ clknet_leaf_40_wb_clk_i _02625_ _00928_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10509_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] net763 net590 vssd1 vssd1
+ vccd1 vccd1 _06773_ sky130_fd_sc_hd__a21o_1
Xhold619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ _04419_ _04428_ _04430_ _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or4_1
X_11489_ _07736_ _07738_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10790__C _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10990__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17069__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16016_ net1377 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14181__B1 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ net2158 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] net821 vssd1 vssd1
+ vccd1 vccd1 _02030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13159_ net2748 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\] net830 vssd1 vssd1
+ vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
XANTENNA__10742__A0 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11176__A1_N net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17967_ clknet_leaf_107_wb_clk_i net1729 _01787_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1308 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13287__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1319 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 net2935
+ sky130_fd_sc_hd__dlygate4sd3_1
X_16918_ clknet_leaf_30_wb_clk_i _02478_ _00781_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11298__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17898_ clknet_leaf_75_wb_clk_i net3189 _01718_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16906__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
X_16849_ clknet_leaf_22_wb_clk_i _02409_ _00712_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09091__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13903__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10030__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09321_ net1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[14\] net872
+ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__A_N team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09252_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\] net850
+ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__and3_1
X_08203_ _04571_ _04575_ _04570_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] net709 net757 vssd1
+ vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_A _07915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08134_ team_01_WB.instance_to_wrap.cpu.f0.state\[5\] team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__nor2_1
XANTENNA__11222__A1 _07256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09828__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11129__A1_N _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12970__A1 _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ team_01_WB.instance_to_wrap.cpu.f0.num\[11\] vssd1 vssd1 vccd1 vccd1 _04496_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1134_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__B _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14172__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout594_A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15565__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1301_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09563__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _05227_ _05228_ _05229_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08898_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\] net739 net693 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\]
+ _05150_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08154__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17831__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14909__A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10860_ _06835_ _07122_ _06777_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09103__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[9\] net718 _05762_ _05765_
+ _05769_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10791_ _06643_ _04935_ net499 vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12530_ net3068 net211 net410 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17981__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12461_ net2917 net309 net418 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14200_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\] _04247_ _04250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\]
+ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__a22o_1
X_11412_ net769 _07441_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09738__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15180_ net1252 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12392_ net2176 net298 net426 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
XANTENNA__11213__B2 _06315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17211__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] _04278_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a22o_1
XANTENNA__12961__A1 net1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ _07020_ _07185_ _07606_ _05014_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09457__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10972__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__B _04624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14163__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nor2_1
X_11274_ _05757_ _06905_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__nand2_1
X_13013_ net2392 net259 net363 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
X_10225_ net1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\] net910 vssd1
+ vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17821_ clknet_leaf_66_wb_clk_i _03378_ _01642_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09473__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] net880 vssd1
+ vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__and3_1
XANTENNA__16929__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13269__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5 _02008_ vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
X_17752_ clknet_leaf_114_wb_clk_i _03310_ _01573_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12103__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ net1021 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] net905 vssd1
+ vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__and3_1
XANTENNA__10412__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14964_ net1243 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08145__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ clknet_leaf_2_wb_clk_i _02263_ _00566_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_13915_ net2669 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[28\]
+ sky130_fd_sc_hd__and2_1
X_17683_ clknet_leaf_74_wb_clk_i _03243_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14895_ net1251 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XANTENNA__11942__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13723__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16634_ clknet_leaf_106_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[20\]
+ _00497_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13846_ _04110_ _04131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08817__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13442__B team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13777_ net1900 net786 _04082_ _04083_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
X_16565_ clknet_leaf_125_wb_clk_i _02193_ _00428_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10989_ _07178_ _07180_ net529 vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ net1280 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12728_ net2986 net210 net386 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16496_ clknet_leaf_106_wb_clk_i _02124_ _00359_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18235_ net1592 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12659_ net2066 net307 net394 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XANTENNA__12773__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15447_ net1243 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11204__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18166_ net1540 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
XFILLER_0_29_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15378_ net1178 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12952__A1 _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17117_ clknet_leaf_128_wb_clk_i _02677_ _00980_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14329_ net2973 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__clkbuf_1
X_18097_ net1471 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__08620__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold416 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold438 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14154__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17048_ clknet_leaf_30_wb_clk_i _02608_ _00911_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold449 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09086__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _06130_ _06131_ _06132_ _06133_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__or4_1
Xfanout907 net909 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_4
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_4
XANTENNA__10025__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout929 net930 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_4
XANTENNA__09581__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\] net731 _05072_
+ _05078_ _05081_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09814__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1116 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08752_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\] net930 vssd1
+ vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__and3_1
Xhold1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12013__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
X_08683_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] net655 net632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08687__A2 _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10494__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\] net753 net735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17234__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\] net752 net717 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12683__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10992__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14464__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_A _03574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1349_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[16\] net962 vssd1
+ vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__and3_1
XANTENNA__09939__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08462__A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14183__B _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08117_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _04500_ team_01_WB.instance_to_wrap.cpu.f0.num\[1\]
+ _04482_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12943__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09097_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] net743 net698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08611__A2 _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14145__B1 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 _04479_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold950 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold961 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[21\] vssd1 vssd1 vccd1 vccd1
+ net2577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ _06270_ _06271_ _06272_ _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__or4_1
XANTENNA__09293__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] net740 _06248_ _06252_
+ _06259_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1650 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 net3266
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11961_ net3141 net313 net473 vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__mux2_1
XANTENNA__12858__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14639__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13671__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] _04021_ vssd1 vssd1 vccd1 vccd1
+ _04022_ sky130_fd_sc_hd__or2_1
X_10912_ net332 _05204_ _05202_ net334 vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14680_ net1405 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XANTENNA__10485__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[1\] net677 net779 vssd1 vssd1
+ vccd1 vccd1 _08003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ _03813_ _03820_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10843_ _06314_ _07084_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__or2_2
XFILLER_0_36_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11063__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16350_ clknet_leaf_65_wb_clk_i net1802 _00218_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
X_13562_ _07903_ _03906_ net185 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10774_ _06485_ _06414_ net505 vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15301_ net1232 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
X_12513_ net2432 net252 net408 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16281_ clknet_leaf_87_wb_clk_i _00012_ _00149_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_18185__1559 vssd1 vssd1 vccd1 vccd1 _18185__1559/HI net1559 sky130_fd_sc_hd__conb_1
XANTENNA__12593__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13493_ _03844_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16601__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18020_ net1597 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09468__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12444_ net3077 net284 net416 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
X_15232_ net1286 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08372__A _04624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15163_ net1298 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12375_ net2303 net200 net423 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XANTENNA__10407__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14136__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14114_ _04224_ _04226_ _04236_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__and3_4
XFILLER_0_107_1643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11326_ _04905_ _06985_ net332 _04906_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__o22ai_1
X_15094_ net1303 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16751__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17877__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14045_ _04213_ net566 _04212_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__and3b_1
XANTENNA__13718__A team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11257_ _07495_ _07510_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_24_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10208_ _06469_ _06470_ _06471_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08311__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ _07450_ _07451_ net541 vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__mux2_1
XANTENNA__17107__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17804_ clknet_leaf_59_wb_clk_i _03361_ _01625_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11238__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] net698 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__a22o_1
X_15996_ net1394 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__inv_2
XANTENNA__08118__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09931__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17735_ clknet_leaf_96_wb_clk_i _03293_ _01556_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14947_ net1219 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XANTENNA__12768__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__A0 _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10476__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17666_ clknet_leaf_144_wb_clk_i _03226_ _01529_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14878_ net1312 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08547__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11673__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17257__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ clknet_leaf_96_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[3\]
+ _00480_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13829_ team_01_WB.instance_to_wrap.cpu.c0.count\[11\] team_01_WB.instance_to_wrap.cpu.c0.count\[8\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] team_01_WB.instance_to_wrap.cpu.c0.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__or4bb_1
XANTENNA__16186__D net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17597_ clknet_leaf_127_wb_clk_i _03157_ _01460_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ clknet_leaf_45_wb_clk_i _02176_ _00411_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13599__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16281__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13900__B net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16479_ clknet_leaf_76_wb_clk_i net2456 _00342_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_09020_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] net926 vssd1
+ vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and3_1
X_18218_ net602 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11701__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09809__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12925__A1 team_01_WB.instance_to_wrap.a1.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18149_ net1523 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12008__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 team_01_WB.instance_to_wrap.a1.ADR_I\[9\] vssd1 vssd1 vccd1 vccd1 net1829
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 team_01_WB.instance_to_wrap.a1.ADR_I\[5\] vssd1 vssd1 vccd1 vccd1 net1851
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 _03328_ vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold257 _01963_ vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _01902_ vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ net987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] net923 vssd1
+ vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout704 net705 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_6
Xfanout726 _04667_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_12
X_09853_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] net938 vssd1
+ vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__and3_1
Xfanout737 _04658_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _04645_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_8
Xfanout759 net762 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
X_08804_ _05067_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__inv_2
XANTENNA__10052__A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\] net723 _04680_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a22o_1
XANTENNA__13102__A1 _06244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08109__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09306__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08735_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\] net660 net616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12678__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14459__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1299_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08666_ _04909_ _04927_ _04928_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11664__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\] net914
+ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16624__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_134_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_hold1574_A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08832__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08904__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ _05448_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09288__A _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[25\] net636 net631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ _05404_ _05410_ _05411_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10927__B1 _07184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12160_ net3159 net300 net450 vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XANTENNA__09793__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08920__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _07311_ _07334_ _07085_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10942__A3 _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ net2457 net314 net456 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
Xhold780 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold791 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11042_ _07300_ _07305_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11352__A0 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15850_ net1198 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14801_ net1361 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15781_ net1229 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12588__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ net2348 net230 net360 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
Xhold1480 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3096 sky130_fd_sc_hd__dlygate4sd3_1
X_17520_ clknet_leaf_23_wb_clk_i _03080_ _01383_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1491 team_01_WB.instance_to_wrap.cpu.K0.code\[2\] vssd1 vssd1 vccd1 vccd1 net3107
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14732_ net1318 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XANTENNA__11655__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11944_ net2621 net223 net473 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17451_ clknet_leaf_60_wb_clk_i _03011_ _01314_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11875_ net2659 net261 net481 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__mux2_1
X_14663_ net1364 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XANTENNA_output107_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16402_ clknet_leaf_102_wb_clk_i net2159 _00265_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10826_ _07088_ _07089_ net516 vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__mux2_1
X_13614_ net188 _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__nand2_1
X_17382_ clknet_leaf_141_wb_clk_i _02942_ _01245_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14594_ net1411 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16333_ clknet_leaf_60_wb_clk_i _01967_ _00201_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13545_ net967 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] _03891_ _03892_
+ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a22o_1
X_10757_ _07011_ _07020_ net538 vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__mux2_1
XANTENNA__09198__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16264_ clknet_leaf_69_wb_clk_i _01901_ _00132_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _03826_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__nor2_1
XANTENNA__08306__S net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10688_ _06861_ _06864_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__or2_2
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09629__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18003_ clknet_leaf_65_wb_clk_i _03552_ _01823_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12907__A1 team_01_WB.instance_to_wrap.a1.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12907__B2 _03608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ net1814 net313 net421 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
XANTENNA__11240__B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15215_ net1246 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16195_ clknet_leaf_87_wb_clk_i _01862_ _00063_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_80_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14109__B1 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13580__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__B1 _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ net2211 net298 net493 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15146_ net1197 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13539__A2_N _07585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11309_ _07070_ _07076_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nor2_1
X_15077_ net1232 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
X_12289_ net3100 net305 net434 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14028_ net3227 net565 _04203_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09000__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09364__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10303__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15979_ net1386 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\] net625 net615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10449__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17718_ clknet_leaf_109_wb_clk_i _03278_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08451_ _04628_ _04635_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__and2_1
X_17649_ clknet_leaf_22_wb_clk_i _03209_ _01512_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08382_ net1120 net956 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__and2_2
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13630__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10746__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_118_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09539__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09003_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[19\] net642 net625 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13020__B1 _07809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout305_A _07970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1047_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13571__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1214_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16177__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13323__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09905_ _06165_ _06166_ _06167_ _06168_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__or4_1
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
Xfanout523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17422__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout534 _06383_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09274__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net547 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11885__A1 _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout567 net569 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_4
X_09836_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\] _04740_ _06088_
+ _06089_ _06091_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__a2111o_1
Xfanout578 net580 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_4
X_18184__1558 vssd1 vssd1 vccd1 vccd1 _18184__1558/HI net1558 sky130_fd_sc_hd__conb_1
Xfanout589 _03585_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09571__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout841_A team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _05963_ _06030_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__or2_1
XANTENNA__17572__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12201__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] net749 net695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a22o_1
X_09698_ _05960_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08649_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[28\] net925 vssd1
+ vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[20\] net1158 net567 net1116
+ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a22o_1
XANTENNA__08915__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ _05166_ _05201_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11591_ _07805_ net496 net2269 net839 vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire902 _04736_ vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_106_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10073__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ net1164 team_01_WB.instance_to_wrap.a1.prev_BUSY_O net798 vssd1 vssd1 vccd1
+ vccd1 _03747_ sky130_fd_sc_hd__and3b_2
X_10542_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ net1749 net816 net600 team_01_WB.instance_to_wrap.a1.ADR_I\[30\] vssd1 vssd1
+ vccd1 vccd1 _02013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[25\] _04650_
+ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15000_ net1256 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
X_12212_ net2629 net285 net441 vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__mux2_1
XANTENNA__09746__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13192_ net3006 net2827 net826 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XANTENNA_input68_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08650__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12143_ net2417 net199 net447 vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13314__A1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09518__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12074_ net2664 net232 net457 vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__mux2_1
X_16951_ clknet_leaf_11_wb_clk_i _02511_ _00814_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11025_ _06607_ _06610_ _05138_ _05206_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__a211o_1
X_15902_ net1346 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__inv_2
XANTENNA__11876__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16882_ clknet_leaf_31_wb_clk_i _02442_ _00745_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10123__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15833_ net1237 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11089__C1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15764_ net1237 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__inv_2
XANTENNA__12111__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12976_ net1832 net605 net587 _03658_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17503_ clknet_leaf_5_wb_clk_i _03063_ _01366_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14715_ net1407 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ net1880 net259 net477 vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ net1251 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XANTENNA__11950__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17434_ clknet_leaf_36_wb_clk_i _02994_ _01297_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14646_ net1375 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
X_11858_ net2332 net315 net480 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10809_ net531 _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__nand2_1
X_17365_ clknet_leaf_8_wb_clk_i _02925_ _01228_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14577_ net1361 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11789_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[20\] net676 net775 vssd1 vssd1
+ vccd1 vccd1 _07919_ sky130_fd_sc_hd__o21a_1
X_16316_ clknet_leaf_81_wb_clk_i _01950_ _00184_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ net767 _07600_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__nor2_1
XANTENNA__11800__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17296_ clknet_leaf_30_wb_clk_i _02856_ _01159_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09359__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16247_ clknet_leaf_86_wb_clk_i _00010_ _00115_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12781__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13459_ _03798_ _03800_ _03803_ _03811_ _03796_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o221a_1
XFILLER_0_109_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09757__B1 _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
X_16178_ clknet_leaf_90_wb_clk_i _01846_ _00046_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
X_15129_ net1238 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08980__A1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10119__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13906__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] net624 _05868_ _05869_
+ _05877_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13069__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09822__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13117__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[9\] net640 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a22o_1
XANTENNA__11619__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08503_ net1003 net907 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__and2_4
XANTENNA__14281__A2 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _05743_ _05744_ _05745_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_1647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout255_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13641__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[31\] net736 _04665_
+ _04673_ _04649_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_52_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08365_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1164_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08799__B2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[60\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09269__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15568__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12691__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13544__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09566__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08470__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16812__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17938__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11307__A0 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1307 net1415 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_4
Xfanout320 _07700_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
Xfanout1318 net1319 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__buf_4
XANTENNA__10224__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1329 net1338 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__clkbuf_4
Xfanout331 _06989_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
Xfanout342 _06979_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_4
Xfanout353 _03751_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout375 _03570_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_8
XFILLER_0_96_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08723__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _03568_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09920__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16962__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout397 _03565_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_6
X_09819_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\] net852 vssd1
+ vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__and3_1
XANTENNA__09732__C _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12830_ net2461 net191 net367 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
XANTENNA__10240__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09279__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14272__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12761_ net2534 net210 net381 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14500_ net1344 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
X_11712_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _07852_ vssd1 vssd1
+ vccd1 vccd1 _07853_ sky130_fd_sc_hd__and2_1
X_12692_ net2883 net308 net390 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15480_ net1255 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08645__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14431_ net1233 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
X_11643_ net1868 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[2\] net841 vssd1 vssd1
+ vccd1 vccd1 _03318_ sky130_fd_sc_hd__mux2_1
XANTENNA__13232__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17150_ clknet_leaf_13_wb_clk_i _02710_ _01013_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11574_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] _07797_ vssd1 vssd1 vccd1 vccd1
+ _07799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14362_ net1382 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17468__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16101_ net1348 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__inv_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
X_13313_ net1704 net810 net805 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\] vssd1
+ vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a22o_1
X_10525_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[24\] net929
+ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__and3_1
X_14293_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\] _04194_ net1804 vssd1
+ vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a21oi_1
X_17081_ clknet_leaf_17_wb_clk_i _02641_ _00944_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13535__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ net50 net39 net64 net61 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__or4_1
X_16032_ net1377 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__inv_2
X_10456_ _06697_ _06718_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12889__A3 _03595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08811__C _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ net2608 net1771 net830 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10387_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\] net654 net647 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__a22o_1
XANTENNA__10415__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12106__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ net2372 net243 net454 vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__mux2_1
X_17983_ clknet_leaf_59_wb_clk_i _03532_ _01803_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11945__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ net2491 net302 net461 vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
X_18032__1426 vssd1 vssd1 vccd1 vccd1 _18032__1426/HI net1426 sky130_fd_sc_hd__conb_1
X_16934_ clknet_leaf_138_wb_clk_i _02494_ _00797_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11008_ _07090_ _07094_ net528 vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16865_ clknet_leaf_138_wb_clk_i _02425_ _00728_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09642__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15816_ net1204 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__inv_2
X_16796_ clknet_leaf_15_wb_clk_i _02356_ _00659_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14263__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15747_ net1220 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12776__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ net1035 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1
+ vccd1 _03646_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13461__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10285__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15678_ net1296 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09690__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17417_ clknet_leaf_41_wb_clk_i _02977_ _01280_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14629_ net1369 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13774__A1 _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ net1660 net550 net347 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1
+ vccd1 vccd1 _03545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17348_ clknet_leaf_128_wb_clk_i _02908_ _01211_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_18183__1557 vssd1 vssd1 vccd1 vccd1 _18183__1557/HI net1557 sky130_fd_sc_hd__conb_1
XANTENNA__09089__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08081_ team_01_WB.instance_to_wrap.cpu.RU0.state\[0\] vssd1 vssd1 vccd1 vccd1 _04510_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17279_ clknet_leaf_2_wb_clk_i _02839_ _01142_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16835__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10028__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09817__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12016__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ net1087 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[19\] net892
+ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout372_A _03571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ net1079 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] net885 vssd1
+ vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__and3_1
XANTENNA__10060__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14254__A2 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] net871 vssd1
+ vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__and3_1
XANTENNA__11068__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12686__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_133_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout637_A _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1379_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\] net910
+ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08465__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17610__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13090__B net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ net973 net920 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__and2_1
XANTENNA__09418__C1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\] net863 vssd1
+ vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08348_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] net2850 net1037 vssd1 vssd1
+ vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XANTENNA__09969__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[69\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10310_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] net932 vssd1
+ vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11290_ net536 _07553_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__nand2_1
X_10241_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\] net859 vssd1
+ vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10172_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\] net862 vssd1
+ vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_100_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1115 net1116 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_1
Xfanout1126 net1140 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_2
XFILLER_0_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1137 net1139 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__buf_2
X_14980_ net1224 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
Xfanout1148 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1
+ net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13931_ net1168 net1058 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[12\] sky130_fd_sc_hd__and3b_1
Xfanout194 net197 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
XANTENNA__09462__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16650_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[4\]
+ _00513_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13862_ team_01_WB.instance_to_wrap.cpu.DM0.dhit team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ _04618_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14245__A2 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15601_ net1192 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XANTENNA__16708__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ net2309 net274 net372 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12596__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16581_ clknet_leaf_65_wb_clk_i _02209_ _00444_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13793_ net1064 _07705_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15532_ net1252 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12744_ net1923 net250 net380 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08375__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15463_ net1183 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
X_12675_ net2086 net282 net387 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17202_ clknet_leaf_31_wb_clk_i _02762_ _01065_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ net1308 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18182_ net1556 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
X_11626_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[13\] _07806_ vssd1 vssd1 vccd1
+ vccd1 _07828_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15394_ net1307 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ clknet_leaf_19_wb_clk_i _02693_ _00996_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1 vssd1 vccd1
+ vccd1 _02253_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07786_ _07787_ vssd1 vssd1 vccd1
+ vccd1 _03357_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08632__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire562 _05052_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13220__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17064_ clknet_leaf_61_wb_clk_i _02624_ _00927_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ _06759_ _06761_ _06771_ net668 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__o32a_4
X_11488_ _07727_ _07734_ net1061 vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__a21o_1
X_14276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[63\] _04253_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[7\]
+ _04158_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09637__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08541__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16015_ net1376 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__inv_2
X_10439_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] net664 net633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[26\]
+ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13227_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] net2383 net825 vssd1 vssd1
+ vccd1 vccd1 _02031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09934__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[76\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10742__A1 _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16238__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12109_ net3191 net287 net451 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
X_13089_ net557 _07807_ _03704_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__o21ai_1
X_17966_ clknet_leaf_98_wb_clk_i _03516_ _01786_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[125\]
+ sky130_fd_sc_hd__dfstp_1
Xhold1309 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16917_ clknet_leaf_26_wb_clk_i _02477_ _00780_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17897_ clknet_leaf_106_wb_clk_i net2062 _01717_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16848_ clknet_leaf_30_wb_clk_i _02408_ _00711_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16388__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14236__A2 _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13903__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16779_ clknet_leaf_46_wb_clk_i _02339_ _00642_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09320_ net1155 net576 net577 vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09251_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] net762 _05513_ _05514_
+ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a22o_4
XFILLER_0_5_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08871__A0 _05133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08202_ net1696 net553 _04568_ _04599_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17783__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ net712 _05438_ _05442_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or4_4
XFILLER_0_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09415__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ _04505_ team_01_WB.instance_to_wrap.cpu.f0.state\[7\] vssd1 vssd1 vccd1 vccd1
+ _04560_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08623__B1 _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout218_A _07943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08064_ team_01_WB.instance_to_wrap.cpu.f0.num\[13\] vssd1 vssd1 vccd1 vccd1 _04495_
+ sky130_fd_sc_hd__inv_2
XANTENNA__10430__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14750__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1127_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout587_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[19\] net685 _05213_
+ _05223_ _05224_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_23_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13683__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout754_A _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] net722 _05141_
+ _05146_ _05149_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10497__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14227__A2 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\] net745 net692 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__a22o_1
X_10790_ net542 net531 _06953_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and3_1
XANTENNA__09654__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] net729 net715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12460_ net2463 net312 net418 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
X_18031__1425 vssd1 vssd1 vccd1 vccd1 _18031__1425/HI net1425 sky130_fd_sc_hd__conb_1
XFILLER_0_47_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11411_ net769 _07669_ net968 vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08614__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ net2087 net244 net425 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14130_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[9\] _04252_ _04280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[97\]
+ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10421__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11342_ _05011_ net336 net333 _07605_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12961__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14061_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__and2b_1
X_11273_ _05755_ _07326_ _05758_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input50_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] net667 vssd1 vssd1
+ vccd1 vccd1 _06488_ sky130_fd_sc_hd__or2_2
X_13012_ net2900 net300 net363 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
X_17820_ clknet_leaf_66_wb_clk_i _03377_ _01641_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_10155_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\] net880 vssd1
+ vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17751_ clknet_leaf_114_wb_clk_i _03309_ _01572_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold6 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 net1622
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] net667 vssd1 vssd1
+ vccd1 vccd1 _06350_ sky130_fd_sc_hd__nor2_1
XANTENNA__09192__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17656__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14963_ net1186 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18182__1556 vssd1 vssd1 vccd1 vccd1 _18182__1556/HI net1556 sky130_fd_sc_hd__conb_1
XFILLER_0_136_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08145__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702_ clknet_leaf_13_wb_clk_i _02262_ _00565_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__B1 _06750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ net2704 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[27\]
+ sky130_fd_sc_hd__and2_1
X_17682_ clknet_leaf_74_wb_clk_i _03242_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14894_ net1222 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
XANTENNA__10131__C _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14218__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16633_ clknet_leaf_105_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[19\]
+ _00496_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13845_ team_01_WB.instance_to_wrap.cpu.c0.count\[1\] team_01_WB.instance_to_wrap.cpu.c0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16564_ clknet_leaf_30_wb_clk_i _02192_ _00427_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13776_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07708_ net782 vssd1 vssd1 vccd1
+ vccd1 _04083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13442__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09645__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10988_ net534 _07251_ _07250_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15515_ net1299 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XANTENNA__08536__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ net2081 net292 net386 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16495_ clknet_leaf_75_wb_clk_i net1768 _00358_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18234_ net603 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15446_ net1260 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ net2362 net311 net394 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18165_ net1539 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_0_111_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11609_ net497 _07819_ net2089 net838 vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__o2bb2a_1
X_15377_ net1199 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
X_12589_ net1921 net243 net401 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__mux2_1
X_17116_ clknet_leaf_15_wb_clk_i _02676_ _00979_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14328_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1
+ vccd1 _02270_ sky130_fd_sc_hd__clkbuf_1
X_18096_ net1470 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold406 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09367__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold417 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\] vssd1 vssd1 vccd1 vccd1
+ net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[4\] vssd1 vssd1 vccd1 vccd1
+ net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15666__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17047_ clknet_leaf_9_wb_clk_i _02607_ _00910_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14259_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\] _04247_ _04266_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[23\]
+ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09664__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_4
Xfanout919 _04675_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_8
X_08820_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\] net727 net715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a22o_1
Xhold1106 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _05013_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__and2_1
Xhold1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ clknet_leaf_106_wb_clk_i _03499_ _01769_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[108\]
+ sky130_fd_sc_hd__dfstp_1
Xhold1139 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\] vssd1 vssd1 vccd1 vccd1
+ net2755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10479__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08682_ _04942_ _04944_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__or3_1
XANTENNA__14209__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13680__A3 _07477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13125__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09097__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ net1130 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\] net922
+ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout335_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1077_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[15\] net936
+ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\] net944 vssd1
+ vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16382__D net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout502_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17529__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1244_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] _04490_ team_01_WB.instance_to_wrap.cpu.f0.num\[23\]
+ _04466_ _04524_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__o221a_1
XANTENNA__14183__C _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09096_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\] net931 vssd1
+ vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08047_ net1065 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14145__B2 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1411_A net1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold940 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold951 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold962 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold973 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold984 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] vssd1 vssd1 vccd1 vccd1
+ net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout871_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout969_A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12204__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[4\] net744 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13656__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ net978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] net924 vssd1
+ vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1
+ net3256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 net3267
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11960_ net2413 net260 net474 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08918__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ _07166_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09740__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net678 _07441_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__nand2_1
X_13630_ net969 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1
+ vccd1 _03964_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11790__A1_N net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _06314_ _07084_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13561_ _03844_ _03905_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10773_ _06485_ net505 vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08835__B1 _05097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14655__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15300_ net1224 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12512_ net2301 net256 net409 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11175__A1_N net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16280_ clknet_leaf_87_wb_clk_i _00011_ _00148_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_137_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13492_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _05064_ vssd1 vssd1
+ vccd1 vccd1 _03845_ sky130_fd_sc_hd__xor2_1
XANTENNA__08653__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ net1293 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ net2825 net222 net417 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08372__B _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15162_ net1265 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
XANTENNA__09187__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12374_ net2391 net288 net423 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
X_14113_ net792 net787 _04232_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__and3_4
XANTENNA__15486__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ net537 _07170_ _07573_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__o21ai_1
X_15093_ net1173 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10126__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14044_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ _04210_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ _07244_ _07511_ _07513_ _07519_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__o211a_2
XFILLER_0_120_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] net751 net739 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12114__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _07387_ _07389_ net529 vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10138_ _06386_ _06400_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__or3_1
X_17803_ clknet_leaf_59_wb_clk_i _03360_ _01624_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_15995_ net1386 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__inv_2
XANTENNA__13647__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13111__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17734_ clknet_leaf_96_wb_clk_i _03292_ _01555_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10069_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[3\] net728 net694 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[3\]
+ _06328_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__a221o_1
X_14946_ net1286 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XANTENNA__11122__A1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17665_ clknet_leaf_135_wb_clk_i _03225_ _01528_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14877_ net1315 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16616_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[2\]
+ _00479_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13828_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04119_ vssd1 vssd1 vccd1
+ vccd1 _04121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17596_ clknet_leaf_11_wb_clk_i _03156_ _01459_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14072__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ clknet_leaf_65_wb_clk_i _02175_ _00410_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13759_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _04015_ _04069_ vssd1 vssd1 vccd1
+ vccd1 _04070_ sky130_fd_sc_hd__o21a_1
XANTENNA__12784__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16426__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16478_ clknet_leaf_85_wb_clk_i net2442 _00341_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18217_ net602 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15429_ net1233 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
XANTENNA__11701__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18148_ net1522 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12925__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16576__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__B1 _05513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[11\] vssd1 vssd1 vccd1 vccd1
+ net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18079_ net1453 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_44_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold225 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold247 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[14\] vssd1 vssd1 vccd1 vccd1
+ net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 net1874
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10036__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold269 team_01_WB.instance_to_wrap.a1.ADR_I\[2\] vssd1 vssd1 vccd1 vccd1 net1885
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _06181_ _06182_ _06183_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__or4_1
XANTENNA__09394__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12689__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 _04681_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_8
XFILLER_0_42_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout716 _04676_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_6
XANTENNA__11429__A team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12024__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[6\] net918 vssd1
+ vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__and3_1
Xfanout727 _04664_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_6
XANTENNA__17971__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 _04643_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_6
X_08803_ _05043_ _05065_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__and2_1
X_09783_ net1143 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[7\] net927 vssd1
+ vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__and3_1
XANTENNA__10052__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18030__1424 vssd1 vssd1 vccd1 vccd1 _18030__1424/HI net1424 sky130_fd_sc_hd__conb_1
XANTENNA_fanout285_A _07920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _04993_ _04995_ _04996_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__or4_1
XANTENNA__11113__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] net746 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout452_A _08018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1194_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08596_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[29\] net963
+ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12694__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13810__B1 _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout717_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09569__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08473__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09217_ _05449_ _05480_ net583 vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08192__B _04592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13574__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18181__1555 vssd1 vssd1 vccd1 vccd1 _18181__1555/HI net1555 sky130_fd_sc_hd__conb_1
XFILLER_0_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09148_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\] net615 _05391_
+ _05399_ _05403_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__B2 _07185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09079_ _05334_ _05335_ _05341_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__or4_2
XFILLER_0_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11110_ _06041_ net341 net337 _05890_ _07373_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__o221a_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net2899 net302 net456 vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold770 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09735__C net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold781 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\] vssd1 vssd1 vccd1 vccd1
+ net2397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11041_ net545 _07295_ _07080_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__o21ba_1
Xhold792 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13341__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11352__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14800_ net1308 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XANTENNA__13554__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15780_ net1272 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__inv_2
X_12992_ net3021 net236 net360 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XANTENNA__08648__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1470 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3097 sky130_fd_sc_hd__dlygate4sd3_1
X_14731_ net1323 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1492 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net3108 sky130_fd_sc_hd__dlygate4sd3_1
X_11943_ net2616 net228 net471 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__mux2_1
XANTENNA__09470__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08367__B net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17450_ clknet_leaf_43_wb_clk_i _03010_ _01313_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08520__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14662_ net1378 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
X_11874_ net778 _07986_ _07987_ _07988_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16401_ clknet_leaf_85_wb_clk_i _02029_ _00264_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13613_ _03814_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__xnor2_1
X_17381_ clknet_leaf_135_wb_clk_i _02941_ _01244_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ _05166_ _05099_ net502 vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__mux2_1
X_14593_ net1403 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16332_ clknet_leaf_63_wb_clk_i net1731 _00200_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13544_ net771 _07152_ net967 vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16599__CLK clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _07014_ _07019_ net530 vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17844__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08814__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16263_ clknet_leaf_69_wb_clk_i _01900_ _00131_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12109__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__inv_2
X_10687_ _04799_ _06947_ _06948_ net323 _06950_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_36_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18002_ clknet_leaf_65_wb_clk_i _03551_ _01822_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_15214_ net1228 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XANTENNA__12907__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ net2272 net259 net422 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16194_ clknet_leaf_87_wb_clk_i _01861_ _00062_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11948__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15145_ net1228 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10819__A_N net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ net2784 net244 net492 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16105__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17994__CLK clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10394__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11591__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ net332 _07570_ _07571_ _06667_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15076_ net1270 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12288_ net2652 net264 net432 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
X_14027_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__or2_1
XANTENNA__13332__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ net535 _07233_ _07502_ _07106_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__o211a_1
XANTENNA__10146__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__A1 _07020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17224__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12779__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13464__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15978_ net1387 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__inv_2
XANTENNA__09839__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17717_ clknet_leaf_109_wb_clk_i _03277_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14929_ net1192 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17374__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] net759 _04712_ _04713_
+ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a22o_1
X_17648_ clknet_leaf_23_wb_clk_i _03208_ _01511_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08381_ net1130 net951 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__and2_4
XFILLER_0_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17579_ clknet_leaf_60_wb_clk_i _03139_ _01442_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11712__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12019__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] net635 _05249_
+ _05251_ _05260_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13020__A1 _06106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13020__B2 _05549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11858__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10385__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08232__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13323__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\] net632 _06151_ _06154_
+ _06161_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11159__A _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout502 net508 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
Xfanout513 _06523_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10063__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout524 _06452_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_2
XANTENNA__10137__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1207_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09852__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] _04745_ _06074_
+ _06079_ _06087_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12689__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout667_A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ _05993_ _06027_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__xnor2_2
XANTENNA__17717__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08717_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\] net731 _04960_
+ _04969_ _04970_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09290__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11637__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09697_ _05923_ _05959_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__or2_1
XANTENNA__10845__A0 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08648_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[28\] net938 vssd1
+ vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__and3_1
XANTENNA__17867__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08579_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] net626 net610 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ _05205_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11590_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\] _07809_ _07808_ vssd1 vssd1
+ vccd1 vccd1 _07810_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10541_ _06796_ _06798_ _06802_ _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__or4_4
XFILLER_0_52_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10238__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16891__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13260_ net1753 net816 net600 team_01_WB.instance_to_wrap.a1.ADR_I\[31\] vssd1 vssd1
+ vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10472_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\] net945
+ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__and3_1
XANTENNA__08569__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11768__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ net2642 net225 net441 vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ net2128 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\] net830 vssd1 vssd1
+ vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__A1 _07702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12142_ net2473 net289 net447 vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09465__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16950_ clknet_leaf_31_wb_clk_i _02510_ _00813_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12073_ net2253 net236 net455 vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__mux2_1
X_15901_ net1346 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__inv_2
X_11024_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__inv_2
X_16881_ clknet_leaf_22_wb_clk_i _02441_ _00744_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13025__A_N net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11876__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12599__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17397__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ net1254 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__inv_2
XANTENNA__08741__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14275__B1 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11089__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__C net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15763_ net1187 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
X_12975_ net365 _03656_ _03657_ net1054 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11008__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14714_ net1411 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17502_ clknet_leaf_4_wb_clk_i _03062_ _01365_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11926_ net2122 net299 net477 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__mux2_1
X_15694_ net1230 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ clknet_leaf_125_wb_clk_i _02993_ _01296_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ net1369 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
X_11857_ _07973_ _07974_ net778 vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__mux2_4
XFILLER_0_129_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11532__A team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10808_ _07060_ _07070_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__or3b_1
X_17364_ clknet_leaf_6_wb_clk_i _02924_ _01227_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14576_ net1366 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XANTENNA__09454__B1 _05716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11788_ net676 _07287_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__nand2_1
X_16315_ clknet_leaf_63_wb_clk_i _01949_ _00183_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08544__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13527_ _07876_ _03877_ net185 vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10739_ _06955_ _06964_ _07000_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__a21o_1
X_17295_ clknet_leaf_124_wb_clk_i _02855_ _01158_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11800__A2 _07243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09937__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16246_ clknet_leaf_86_wb_clk_i _00009_ _00114_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13002__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ _03805_ _03807_ _03804_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08841__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ net2448 net228 net419 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16177_ clknet_leaf_90_wb_clk_i _01845_ _00045_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_109_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13389_ team_01_WB.instance_to_wrap.cpu.f0.num\[9\] net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__10367__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15128_ net1259 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15059_ net1188 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XANTENNA__16614__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__A2 _06381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09672__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13906__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11707__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\] net656 _05863_ _05870_
+ _05871_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08732__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__A1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14266__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16764__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _05811_ _05812_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nor4_1
X_18180__1554 vssd1 vssd1 vccd1 vccd1 _18180__1554/HI net1554 sky130_fd_sc_hd__conb_1
X_08502_ net1002 net881 vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and2_4
XFILLER_0_91_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14281__A3 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09482_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[12\] net653 _05725_
+ _05727_ _05736_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08433_ net984 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[31\] net927 vssd1
+ vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10757__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08364_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\] vssd1 vssd1 vccd1 vccd1 _04628_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10058__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[61\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout415_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09847__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11004__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1324_A net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__B net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08971__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout310 _07998_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11307__A1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1308 net1310 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__buf_4
Xfanout1319 net1325 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout321 _06954_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_4
Xfanout332 _06989_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
Xfanout343 _06979_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 net355 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
Xfanout365 _03582_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 _03570_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_4
XANTENNA__08723__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout387 _03567_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
X_09818_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\] net862 vssd1
+ vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout398 _03565_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_4
XANTENNA__10521__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14257__B1 _04412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10530__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09749_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[10\] net648 net612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a22o_1
XANTENNA__12807__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ net2493 net292 net381 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11711_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ _07851_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12691_ net1962 net313 net390 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14430_ net1233 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
X_11642_ net2107 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] net841 vssd1 vssd1
+ vccd1 vccd1 _03319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ net1382 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
X_11573_ _07702_ _07797_ net320 vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14663__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16100_ net1403 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__inv_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13312_ net1872 net809 net803 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\] vssd1
+ vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
X_17080_ clknet_leaf_27_wb_clk_i _02640_ _00943_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10524_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[24\] net940
+ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14292_ _04201_ _04440_ net1367 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16031_ net1376 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__inv_2
X_13243_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13535__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10455_ _06697_ _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13174_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[60\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09195__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10386_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\] net663 net619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[27\]
+ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08962__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ net3028 net314 net453 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17982_ clknet_leaf_57_wb_clk_i _03531_ _01802_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10134__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12056_ net2822 net264 net461 vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
X_16933_ clknet_leaf_131_wb_clk_i _02493_ _00796_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09923__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09911__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13218__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _06970_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__and2_1
XANTENNA__12122__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16864_ clknet_leaf_2_wb_clk_i _02424_ _00727_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14248__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08539__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15815_ net1180 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__inv_2
X_16795_ clknet_leaf_39_wb_clk_i _02355_ _00658_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11961__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15746_ net1267 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
X_12958_ net1033 _07368_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__nand2_1
XANTENNA__13471__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ net3001 net200 net475 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
X_15677_ net1284 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12889_ net366 _03594_ _03595_ net1056 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\]
+ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17416_ clknet_leaf_45_wb_clk_i _02976_ _01279_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14628_ net1399 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17412__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17347_ clknet_leaf_133_wb_clk_i _02907_ _01210_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12792__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ net1409 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
XANTENNA__10309__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[3\] vssd1 vssd1 vccd1 vccd1
+ _04509_ sky130_fd_sc_hd__inv_2
XANTENNA__12982__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17278_ clknet_leaf_12_wb_clk_i _02838_ _01141_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16229_ clknet_leaf_38_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[10\]
+ _00097_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08982_ net1085 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\] net863
+ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13128__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12032__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14239__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[8\] net857 vssd1
+ vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14748__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09534_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\] net860 vssd1
+ vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09465_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] net885 vssd1
+ vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1274_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__B net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08416_ net1121 net935 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__and2_4
XFILLER_0_4_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17092__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] net877
+ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08347_ net2731 net2298 net1048 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
XANTENNA__13765__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17905__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08641__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08278_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] net2130 net1040 vssd1 vssd1
+ vccd1 vccd1 _03469_ sky130_fd_sc_hd__mux2_1
XANTENNA__08481__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08912__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12207__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10516__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10240_ net1006 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[1\] net864 vssd1
+ vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__and3_1
XANTENNA__14190__A2 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[2\] net906 vssd1
+ vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1
+ net1105 sky130_fd_sc_hd__clkbuf_8
Xfanout1116 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[20\] vssd1 vssd1 vccd1 vccd1
+ net1116 sky130_fd_sc_hd__clkbuf_4
Xfanout1127 net1140 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09743__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_2
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13930_ net1167 net1060 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[11\] sky130_fd_sc_hd__and3b_1
XFILLER_0_22_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10503__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 net197 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlymetal6s2s_1
X_13861_ _04119_ _04138_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15600_ net1250 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
X_12812_ net2518 net218 net371 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16580_ clknet_leaf_57_wb_clk_i _02208_ _00443_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ net1064 _07705_ net484 vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17435__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15531_ net1206 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
X_12743_ net3124 net255 net379 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08375__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15462_ net1274 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
X_12674_ net2450 net224 net389 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
XANTENNA__09409__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17201_ clknet_leaf_24_wb_clk_i _02761_ _01064_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14413_ net1308 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
X_18181_ net1555 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ net1863 net839 _07808_ _07827_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15393_ net1288 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10129__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ clknet_leaf_47_wb_clk_i _02692_ _00995_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12964__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] vssd1 vssd1 vccd1
+ vccd1 _02254_ sky130_fd_sc_hd__clkbuf_1
X_11556_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _07732_ _07785_ vssd1 vssd1 vccd1
+ vccd1 _07787_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire574 _06380_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
XANTENNA__14166__C1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10507_ _06765_ _06767_ _06769_ _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__or4_1
X_17063_ clknet_leaf_126_wb_clk_i _02623_ _00926_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12117__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14275_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\] _04260_ _04276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[47\]
+ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a221o_1
X_11487_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] _07736_ _07737_ vssd1 vssd1 vccd1
+ vccd1 _03377_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_111_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10990__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16014_ net1358 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__inv_2
X_13226_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[8\] net2164 net823 vssd1 vssd1
+ vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
X_10438_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] net637 net612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11956__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[77\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
X_10369_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[27\] net728 _06617_
+ _06622_ _06625_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16113__A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ net3127 net230 net451 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
X_13088_ net355 _03711_ _03712_ net835 net2693 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a32o_1
X_17965_ clknet_leaf_106_wb_clk_i _03515_ _01785_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[124\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11257__A _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ net3086 net202 net460 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
X_16916_ clknet_leaf_9_wb_clk_i _02476_ _00779_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17896_ clknet_leaf_101_wb_clk_i net1766 _01716_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12787__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16847_ clknet_leaf_124_wb_clk_i _02407_ _00710_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16778_ clknet_leaf_43_wb_clk_i _02338_ _00641_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10258__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15729_ net1199 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XANTENNA__11704__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17928__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] net710 net758 vssd1
+ vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08201_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _04598_ _04567_ vssd1 vssd1 vccd1
+ vccd1 _04599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09181_ _05432_ _05433_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11720__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ net1764 net785 _04559_ team_01_WB.instance_to_wrap.cpu.f0.i\[0\] vssd1 vssd1
+ vccd1 vccd1 _03559_ sky130_fd_sc_hd__a22o_1
XANTENNA__09397__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09828__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16952__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ team_01_WB.instance_to_wrap.cpu.f0.num\[16\] vssd1 vssd1 vccd1 vccd1 _04494_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12027__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09179__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14172__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09033__D1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17308__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1022_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] net749 _05216_
+ _05218_ _05221_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08240__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08896_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\] net740 net736 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17458__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1391_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08476__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] net715 net700 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08907__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout914_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09448_ _05693_ _05709_ _05710_ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09379_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] net746 _05625_
+ _05626_ _05631_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11410_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] _06526_ _07673_ vssd1
+ vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12390_ net2667 net314 net424 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XANTENNA__09738__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14148__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ net339 net342 _05013_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10972__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14060_ net3122 _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__o21a_1
XANTENNA__14163__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11272_ _05755_ _05758_ _07326_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13011_ net2316 net244 net361 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10223_ net781 _04715_ net681 net1113 vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o31a_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input43_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10154_ net1017 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[2\] net909 vssd1
+ vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09473__C net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11077__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17750_ clknet_leaf_114_wb_clk_i _03308_ _01571_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14962_ net1174 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
Xhold7 team_01_WB.instance_to_wrap.a1.ADR_I\[6\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net581 _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__or2_1
XANTENNA__10412__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ clknet_leaf_123_wb_clk_i _02261_ _00564_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13913_ net2923 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[26\]
+ sky130_fd_sc_hd__and2_1
X_17681_ clknet_leaf_74_wb_clk_i _03241_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14893_ net1222 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XANTENNA__08550__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13844_ net2050 _04110_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[2\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12400__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16632_ clknet_leaf_105_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[18\]
+ _00495_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08817__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ net484 _07710_ _04081_ net563 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16563_ clknet_leaf_11_wb_clk_i _02191_ _00426_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ _07164_ _07172_ net526 vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__mux2_1
XANTENNA__11988__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12726_ net2561 net296 net386 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15514_ net1259 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16494_ clknet_leaf_80_wb_clk_i net1641 _00357_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16975__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18233_ net1591 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
X_15445_ net1176 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ net2116 net260 net393 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12937__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[22\] net572 vssd1 vssd1 vccd1
+ vccd1 _07819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18164_ net1538 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_0_136_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15376_ net1262 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
X_12588_ net2228 net314 net400 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08325__S net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17115_ clknet_leaf_39_wb_clk_i _02675_ _00978_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14327_ net1645 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16205__CLK clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15947__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18095_ net1469 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
X_11539_ net1065 _07705_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__nand2_2
Xhold407 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold418 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\] vssd1 vssd1 vccd1 vccd1
+ net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17046_ clknet_leaf_30_wb_clk_i _02606_ _00909_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14154__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14258_ net790 net788 net787 _04393_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a31o_1
Xhold429 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13209_ net3176 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] net829 vssd1 vssd1
+ vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13467__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13362__B1 _03747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\] _04238_ _04255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\]
+ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout909 _04731_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16355__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17600__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15682__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1107 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ _04988_ _05011_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__or2_1
X_17948_ clknet_leaf_81_wb_clk_i net2481 _01768_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[107\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13665__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09680__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08681_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\] net634 net619 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\]
+ _04936_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17879_ clknet_leaf_102_wb_clk_i _03429_ _01699_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11715__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09302_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] net951 vssd1
+ vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\] net917 vssd1
+ vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_A _07897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13141__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\] net922 vssd1
+ vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08235__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08115_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] _04497_ team_01_WB.instance_to_wrap.cpu.f0.num\[3\]
+ _04481_ _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17130__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10066__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09095_ net1127 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\] net963
+ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1237_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08046_ team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 _04477_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09855__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold930 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[72\] vssd1 vssd1 vccd1 vccd1
+ net2546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout697_A _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold952 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] vssd1 vssd1 vccd1 vccd1
+ net2568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13353__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold963 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1404_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold985 _03477_ vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09572__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17280__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\] net926 vssd1
+ vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__and3_1
XANTENNA__09293__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13105__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16848__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _05207_ _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1630 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3246 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09590__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1641 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11667__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1652 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net3268
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08879_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[21\] net938 vssd1
+ vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10910_ net533 _07173_ _06995_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12220__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ net1936 net294 net480 vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ net522 _07104_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14936__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13560_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _05064_ _03904_ vssd1
+ vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08835__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ _07034_ _07035_ net517 vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__mux2_1
X_12511_ net2364 net219 net409 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ _03842_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ net1297 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XANTENNA__12919__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ net2215 net228 net415 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09468__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15161_ net1192 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12373_ net2958 net232 net425 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XANTENNA__14671__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10407__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10945__A2 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\] _04272_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14136__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09765__A _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ _06942_ _06944_ _06840_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__and3b_1
X_15092_ net1240 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13344__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14043_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04210_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__a21o_1
X_11255_ _07517_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10206_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] net743 _06459_ _06461_
+ _06463_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _07386_ _07449_ net523 vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17802_ clknet_leaf_59_wb_clk_i _03359_ _01623_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_10137_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] net688 _06389_ _06390_
+ _06398_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13647__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15994_ net1388 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__inv_2
XANTENNA__09315__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11658__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17733_ clknet_leaf_98_wb_clk_i _03291_ _01554_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_10068_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[3\] net716 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a22o_1
X_14945_ net1312 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09931__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__A2 _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13226__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17664_ clknet_leaf_2_wb_clk_i _03224_ _01527_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ net1315 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08547__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16615_ clknet_leaf_97_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[1\]
+ _00478_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13827_ team_01_WB.instance_to_wrap.cpu.c0.count\[15\] _04119_ vssd1 vssd1 vccd1
+ vccd1 _04120_ sky130_fd_sc_hd__or2_1
X_17595_ clknet_leaf_35_wb_clk_i _03155_ _01458_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16546_ clknet_leaf_64_wb_clk_i _02174_ _00409_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13758_ _07716_ _07773_ _04558_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08844__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12709_ net2007 net221 net383 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16477_ clknet_leaf_79_wb_clk_i _02105_ _00340_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_13689_ _04011_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18216_ net601 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15428_ net1270 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12386__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18147_ net1521 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
X_15359_ net1297 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
XANTENNA__15677__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09251__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09675__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold204 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[7\] vssd1 vssd1 vccd1 vccd1
+ net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\] vssd1 vssd1 vccd1 vccd1
+ net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18078_ net1452 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_123_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold226 net91 vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold237 net75 vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold248 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[4\] vssd1 vssd1 vccd1 vccd1
+ net1864 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\] net740 net732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a22o_1
XANTENNA__13335__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold259 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ clknet_leaf_131_wb_clk_i _02589_ _00892_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12305__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 _04680_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_8
XFILLER_0_106_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[6\] net931 vssd1
+ vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__and3_1
XANTENNA__09554__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 _04674_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_8
Xfanout728 _04664_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _04656_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_8
X_08802_ _05043_ _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__nor2_1
X_09782_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\] net918 vssd1
+ vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09306__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11649__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\] net650 net648 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a22o_1
XANTENNA__08514__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13136__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12040__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[28\] net747 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a22o_1
XANTENNA__10321__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] _04650_
+ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout445_A _08020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1187_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout612_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08473__B net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ _05476_ _05478_ _05479_ _05450_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__o31a_4
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16520__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09147_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] net627 _05384_ _05386_
+ _05394_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_126_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10388__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10227__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09078_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[18\] net640 _05314_ _05318_
+ _05320_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09793__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout981_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13326__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08920__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16670__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12215__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17796__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold760 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\] vssd1 vssd1 vccd1 vccd1
+ net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _05069_ _06876_ _07159_ _07303_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__o31a_1
Xhold793 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11818__A1_N net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13629__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10560__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12991_ net3142 net204 net361 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
Xhold1460 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\] vssd1 vssd1 vccd1 vccd1
+ net3076 sky130_fd_sc_hd__dlygate4sd3_1
X_14730_ net1318 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1471 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3087 sky130_fd_sc_hd__dlygate4sd3_1
X_11942_ net2214 net199 net471 vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__mux2_1
Xhold1482 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net3109 sky130_fd_sc_hd__dlygate4sd3_1
X_14661_ net1369 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
X_11873_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\] net677 net778 vssd1 vssd1
+ vccd1 vccd1 _07988_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17176__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16400_ clknet_leaf_104_wb_clk_i _02028_ _00263_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_13612_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\] _05584_ _03948_ vssd1
+ vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10824_ _04988_ _05043_ net500 vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__mux2_1
X_14592_ net1407 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
X_17380_ clknet_leaf_138_wb_clk_i _02940_ _01243_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16331_ clknet_leaf_63_wb_clk_i net1860 _00199_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
X_13543_ net185 _03889_ _03890_ net771 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a211o_1
X_10755_ _07016_ _07018_ net511 vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__mux2_2
XFILLER_0_137_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16262_ clknet_leaf_71_wb_clk_i _01899_ _00130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_18149__1523 vssd1 vssd1 vccd1 vccd1 _18149__1523/HI net1523 sky130_fd_sc_hd__conb_1
XFILLER_0_129_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13474_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _05449_ vssd1 vssd1
+ vccd1 vccd1 _03827_ sky130_fd_sc_hd__xor2_1
XANTENNA__09198__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ _06947_ _06948_ _04799_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13565__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18001_ clknet_leaf_65_wb_clk_i _03550_ _01821_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15213_ net1212 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12425_ net2757 net298 net422 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
X_16193_ clknet_leaf_92_wb_clk_i _01860_ _00061_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14109__A2 _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09495__A _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144_ net1183 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
X_12356_ net2849 net316 net490 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09784__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13317__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ net338 net340 _06665_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__mux2_1
X_15075_ net1223 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
X_12287_ net3105 net266 net434 vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XANTENNA__12125__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14026_ net3256 net565 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__and2b_1
X_11238_ net541 _07451_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__or2_1
XANTENNA__11964__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__A2 _07185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11169_ _06881_ _07431_ _07432_ net345 vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10551__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18105__1479 vssd1 vssd1 vccd1 vccd1 _18105__1479/HI net1479 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09661__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15977_ net1386 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ clknet_leaf_109_wb_clk_i _03276_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11049__A2_N net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14928_ net1262 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17647_ clknet_leaf_124_wb_clk_i _03207_ _01510_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14859_ net1341 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13480__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08380_ net1149 net1151 net1153 net1147 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_50_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17578_ clknet_leaf_41_wb_clk_i _03138_ _01441_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17669__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16529_ clknet_leaf_59_wb_clk_i _02157_ _00392_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08680__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\] net638 net626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13020__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15200__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13308__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12035__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17049__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[6\] net645 _06148_ _06149_
+ _06153_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11159__B _06867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net508 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_4
Xfanout514 net519 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout525 net527 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_4
Xfanout536 _06383_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08735__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _06314_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_127_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09834_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[7\] net621 _06077_ _06083_
+ _06094_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1102_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08749__A _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 _07836_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_2
X_09765_ _05993_ _06027_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09571__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08468__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15870__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08716_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\] net745 _04964_ _04966_
+ _04968_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_55_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09696_ _05923_ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10845__A1 _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08647_ net1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\] net923
+ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout827_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08578_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] net635 _04840_
+ _04841_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08915__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13795__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10519__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10073__A2 _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[24\] net701 _06779_ _06803_
+ net711 vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11270__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13547__B1 _07669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10471_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[25\] net914
+ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12210_ net2229 net227 net439 vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__mux2_1
X_13190_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[44\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[52\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09746__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08650__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net3179 net232 net449 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__mux2_1
XANTENNA__10781__A0 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09518__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ net2514 net202 net457 vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
Xhold590 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12522__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _07154_ _07266_ _07284_ _07286_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__o211a_4
XFILLER_0_25_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15900_ net1348 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16880_ clknet_leaf_24_wb_clk_i _02440_ _00743_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10533__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15831_ net1238 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15780__A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12974_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[3\] net1035 vssd1 vssd1 vccd1
+ vccd1 _03657_ sky130_fd_sc_hd__or2_1
X_15762_ net1174 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
XANTENNA__16566__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18047__1609 vssd1 vssd1 vccd1 vccd1 net1609 _18047__1609/LO sky130_fd_sc_hd__conb_1
Xhold1290 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ clknet_leaf_127_wb_clk_i _03061_ _01364_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14713_ net1408 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XANTENNA__17811__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ net2999 net244 net478 vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__mux2_1
X_15693_ net1218 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17432_ clknet_leaf_30_wb_clk_i _02992_ _01295_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14644_ net1373 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[8\] _07379_ net677 vssd1 vssd1
+ vccd1 vccd1 _07974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08394__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13786__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ net549 net509 vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__nand2_1
X_17363_ clknet_leaf_49_wb_clk_i _02923_ _01226_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14575_ net1362 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11787_ _07859_ _07916_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__or2_1
XANTENNA__09454__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16314_ clknet_leaf_112_wb_clk_i _01948_ _00182_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13526_ _03865_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17961__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ net542 _06995_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__nand2_1
X_17294_ clknet_leaf_52_wb_clk_i _02854_ _01157_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11959__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13538__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16245_ clknet_leaf_86_wb_clk_i _00008_ _00113_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_13457_ _03803_ _03806_ _03809_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__or3_1
X_10669_ _06919_ _06929_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16116__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12408_ net2978 net198 net419 vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XANTENNA__09757__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ net2697 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1
+ vccd1 vccd1 _01895_ sky130_fd_sc_hd__a22o_1
X_16176_ clknet_leaf_91_wb_clk_i _01844_ _00044_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
X_12339_ net3072 net233 net492 vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
X_15127_ net1244 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__09509__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15058_ net1180 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XANTENNA__09953__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14009_ net160 net71 net73 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__and3b_1
XFILLER_0_78_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17341__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11707__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16909__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[9\] net648 _05801_ _05803_
+ _05807_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a2111o_1
X_18059__1435 vssd1 vssd1 vccd1 vccd1 _18059__1435/HI net1435 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08501_ net1084 net872 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__and2_4
XFILLER_0_37_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09481_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[12\] net628 _05728_
+ _05729_ _05735_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_91_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11723__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ net982 net927 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__and2_4
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] net781 vssd1 vssd1 vccd1
+ vccd1 _04627_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ net2198 net2647 net1040 vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11869__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout310_A _07998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1052_A team_01_WB.instance_to_wrap.cpu.SR1.enable vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08243__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10763__A0 _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1309 net1310 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__buf_2
XANTENNA__08708__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net325 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout333 _06988_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10515__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_4
Xfanout366 _03582_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09920__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 _03570_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_8
X_09817_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[7\] net884 vssd1
+ vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__and3_1
Xfanout388 _03567_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17834__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18148__1522 vssd1 vssd1 vccd1 vccd1 _18148__1522/HI net1522 sky130_fd_sc_hd__conb_1
XFILLER_0_96_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout944_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _03564_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_8
XFILLER_0_119_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09748_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[10\] net891
+ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10240__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10818__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09679_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] net894
+ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11710_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _07850_ vssd1 vssd1 vccd1
+ vccd1 _07851_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12690_ net2989 net260 net389 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08645__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13768__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ net1864 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[4\] net841 vssd1 vssd1
+ vccd1 vccd1 _03320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ net1382 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
XANTENNA__11243__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\] _07795_ vssd1 vssd1 vccd1 vccd1
+ _07797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17214__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ net1725 net808 net804 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[13\] vssd1
+ vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10523_ net971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[24\] net920 vssd1
+ vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__and3_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_14291_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[4\] _04194_ vssd1 vssd1 vccd1
+ vccd1 _04440_ sky130_fd_sc_hd__xnor2_1
X_18104__1478 vssd1 vssd1 vccd1 vccd1 _18104__1478/HI net1478 sky130_fd_sc_hd__conb_1
XFILLER_0_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13242_ _03726_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\] net828 vssd1 vssd1
+ vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
X_16030_ net1358 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__inv_2
XANTENNA_input73_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _06716_ _06717_ net578 vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[61\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10385_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\] net661 net641 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ net2974 net304 net453 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux2_1
XANTENNA__10415__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17981_ clknet_leaf_59_wb_clk_i _03530_ _01801_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12055_ net1990 net267 net462 vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
X_16932_ clknet_leaf_129_wb_clk_i _02492_ _00795_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12403__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _07104_ _07269_ net522 vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__mux2_1
X_18040__1430 vssd1 vssd1 vccd1 vccd1 _18040__1430/HI net1430 sky130_fd_sc_hd__conb_1
XANTENNA__09911__A2 _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16863_ clknet_leaf_5_wb_clk_i _02423_ _00726_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15814_ net1271 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__inv_2
X_16794_ clknet_leaf_33_wb_clk_i _02354_ _00657_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15745_ net1290 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12957_ net1642 net606 net588 _03644_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13234__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10285__A2 _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11908_ net3055 net286 net475 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15676_ net1279 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12888_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] vssd1 vssd1 vccd1
+ vccd1 _03595_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17415_ clknet_leaf_120_wb_clk_i _02975_ _01278_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14627_ net1347 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
X_11839_ net678 _07568_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09978__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17346_ clknet_leaf_143_wb_clk_i _02906_ _01209_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14558_ net1399 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
XANTENNA__08635__C1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13509_ _03760_ _03761_ _03860_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__or3b_1
X_17277_ clknet_leaf_128_wb_clk_i _02837_ _01140_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14489_ net1399 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XANTENNA__10993__B1 _07256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16228_ clknet_leaf_38_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[9\]
+ _00096_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12734__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ clknet_leaf_90_wb_clk_i _01827_ _00027_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10745__A0 _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09683__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[19\] net669 vssd1 vssd1
+ vccd1 vccd1 _05245_ sky130_fd_sc_hd__or2_1
XANTENNA__16731__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17857__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11718__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08166__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09902__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11170__A0 _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09602_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[8\] net860 vssd1
+ vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16881__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10060__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09533_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\] net863 vssd1
+ vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout260_A _07989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13144__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11453__A team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\] net860
+ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17237__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ net985 _04677_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09395_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\] net845
+ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1267_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[10\] net3151 net1048 vssd1 vssd1
+ vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux2_1
XANTENNA__09858__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08762__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16261__CLK clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ net2873 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\] net1045 vssd1 vssd1
+ vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XANTENNA__08641__A2 _04902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__A0 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08481__B net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14175__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09296__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_142_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_18046__1608 vssd1 vssd1 vccd1 vccd1 net1608 _18046__1608/LO sky130_fd_sc_hd__conb_1
XFILLER_0_123_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10235__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] net887 vssd1
+ vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_2
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12223__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1128 net1140 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_2
Xfanout1139 net1140 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_2
XANTENNA__08157__B2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net197 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13860_ net3265 _04118_ net1963 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__a21oi_1
X_12811_ net2690 net279 net372 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ net1686 net782 _04092_ _04094_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ net1198 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
X_12742_ net2971 net221 net379 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15461_ net1232 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
X_12673_ net2593 net226 net387 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17200_ clknet_leaf_24_wb_clk_i _02760_ _01063_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14412_ net1310 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
X_11624_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[14\] _07806_ vssd1 vssd1 vccd1
+ vccd1 _07827_ sky130_fd_sc_hd__and2_1
X_18180_ net1554 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
XFILLER_0_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15392_ net1251 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ clknet_leaf_56_wb_clk_i _02691_ _00994_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12964__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11555_ net483 _07785_ net319 vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__a21o_1
XANTENNA__12964__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14343_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1
+ vccd1 _02255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08632__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10707__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\] _04745_ net629
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[25\] _06754_ vssd1 vssd1 vccd1
+ vccd1 _06770_ sky130_fd_sc_hd__a221o_1
X_17062_ clknet_leaf_139_wb_clk_i _02622_ _00925_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_18058__1434 vssd1 vssd1 vccd1 vccd1 _18058__1434/HI net1434 sky130_fd_sc_hd__conb_1
X_14274_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[39\] _04238_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\]
+ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a22o_1
X_11486_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] _07728_ _07732_ vssd1 vssd1 vccd1
+ vccd1 _07737_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire575 _05684_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_1
XANTENNA__16754__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11519__A2 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13225_ net1720 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] net829 vssd1 vssd1
+ vccd1 vccd1 _02033_ sky130_fd_sc_hd__mux2_1
X_16013_ net1355 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10437_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[26\] net631 net626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\]
+ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ net2718 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\] net820 vssd1 vssd1
+ vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\] net719 net713 vssd1
+ vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09934__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ net2878 net236 net451 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XANTENNA__13229__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12133__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[11\] net1029 vssd1 vssd1 vccd1
+ vccd1 _03712_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17964_ clknet_leaf_81_wb_clk_i net1722 _01784_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10299_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[0\] _04666_ vssd1
+ vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__and3_1
XANTENNA__08148__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16915_ clknet_leaf_49_wb_clk_i _02475_ _00778_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12038_ net3117 net238 net459 vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
XANTENNA__11257__B _07510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17895_ clknet_leaf_107_wb_clk_i _03445_ _01715_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11152__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11972__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13753__A team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16846_ clknet_leaf_55_wb_clk_i _02406_ _00709_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16777_ clknet_leaf_38_wb_clk_i _02337_ _00640_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _04171_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10258__A2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15728_ net1250 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15659_ net1208 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14584__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08200_ _04574_ _04582_ _04585_ _04589_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__or4_2
XFILLER_0_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09678__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] net701 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08131_ net1810 net785 _04559_ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] vssd1 vssd1
+ vccd1 vccd1 _03560_ sky130_fd_sc_hd__a22o_1
XANTENNA__12955__A1 _07379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17329_ clknet_leaf_20_wb_clk_i _02889_ _01192_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12308__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08623__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18147__1521 vssd1 vssd1 vccd1 vccd1 _18147__1521/HI net1521 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14157__B1 _04276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08062_ team_01_WB.instance_to_wrap.cpu.f0.num\[20\] vssd1 vssd1 vccd1 vccd1 _04493_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_113_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10430__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13380__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12043__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[19\] net726 _05215_
+ _05217_ _05220_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10352__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1015_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08895_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[21\] net747 net743 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a22o_1
XANTENNA__11143__A0 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout475_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10497__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103__1477 vssd1 vssd1 vccd1 vccd1 _18103__1477/HI net1477 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08757__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout642_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08476__B net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16627__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[9\] net731 _05764_ _05767_
+ _05772_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\] net752 _05695_ _05697_
+ _05699_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08862__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] net739 net691 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\] net1917 net1051 vssd1 vssd1
+ vccd1 vccd1 _03418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11630__B _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12218__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08614__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ _06877_ _07303_ _07603_ _05015_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10421__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10709__A0 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ net345 _07204_ _07523_ _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__o31a_2
X_13010_ net3087 net317 net362 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10222_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] net765 vssd1 vssd1 vccd1 vccd1
+ _06486_ sky130_fd_sc_hd__and2_1
XANTENNA__13371__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_105_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10153_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] net894 vssd1
+ vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13950__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17402__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ net1200 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
X_10084_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] net765 _04723_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__a22o_1
Xhold8 _01989_ vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13573__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16700_ clknet_leaf_14_wb_clk_i _02260_ _00563_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13912_ net2558 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[25\]
+ sky130_fd_sc_hd__and2_1
X_17680_ clknet_leaf_74_wb_clk_i _03240_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10488__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12882__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ net1307 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16631_ clknet_leaf_116_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[17\]
+ _00494_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13843_ _04111_ _04130_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[3\]
+ sky130_fd_sc_hd__and2b_1
XANTENNA__11805__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11437__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17552__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ clknet_leaf_32_wb_clk_i _02190_ _00425_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13774_ _04472_ _07774_ _04014_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a21oi_1
X_10986_ net539 _07249_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15513_ net1193 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
X_12725_ net3254 net309 net386 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ clknet_leaf_78_wb_clk_i net1634 _00356_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12917__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18232_ net602 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09498__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15444_ net1241 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XANTENNA__13330__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ net2100 net299 net394 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__C _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18163_ net1537 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
X_11607_ net496 _07818_ net2083 net838 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12128__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ net2564 net302 net400 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
X_15375_ net1251 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XANTENNA__08605__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17114_ clknet_leaf_32_wb_clk_i _02674_ _00977_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14139__B1 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14326_ _04169_ _04187_ _04189_ _04167_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11538_ _04475_ _07772_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__nor2_2
X_18094_ net1468 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold408 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ clknet_leaf_26_wb_clk_i _02605_ _00908_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold419 _02143_ vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\] team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ team_01_WB.instance_to_wrap.cpu.f0.i\[1\] team_01_WB.instance_to_wrap.cpu.f0.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14257_ net1706 net585 _04412_ net1171 vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13362__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ net2178 net1646 net826 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09030__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14188_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\] _04227_ _04288_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__a22o_1
XANTENNA__15963__A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ net1663 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\] net824 vssd1 vssd1
+ vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09961__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
X_17947_ clknet_leaf_85_wb_clk_i net1799 _01767_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11125__A0 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12798__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1119 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[96\] vssd1 vssd1 vccd1 vccd1
+ net2735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10479__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[28\] net628 _04943_
+ net670 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__a211o_1
XANTENNA__12873__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17878_ clknet_leaf_98_wb_clk_i _03428_ _01698_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[37\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16829_ clknet_leaf_127_wb_clk_i _02389_ _00692_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11715__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18045__1607 vssd1 vssd1 vccd1 vccd1 net1607 _18045__1607/LO sky130_fd_sc_hd__conb_1
XFILLER_0_53_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09097__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[14\] net930 vssd1
+ vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__and3_1
XANTENNA__13930__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ net973 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[15\] net921 vssd1
+ vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11450__B team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09163_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] net944
+ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__and3_1
XANTENNA__12928__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13050__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_A _07915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08114_ _04478_ team_01_WB.instance_to_wrap.cpu.f0.num\[7\] _04499_ team_01_WB.instance_to_wrap.cpu.f0.i\[3\]
+ _04530_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[17\] net942
+ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08045_ team_01_WB.instance_to_wrap.cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _04476_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold920 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold931 _03471_ vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13353__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold942 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net2558
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold953 _02038_ vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17425__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold964 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold986 team_01_WB.instance_to_wrap.cpu.f0.num\[0\] vssd1 vssd1 vccd1 vccd1 net2602
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09996_ net991 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[4\] net922 vssd1
+ vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__and3_1
XANTENNA__09309__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _05070_ _05210_ _05209_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout857_A _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1642 team_01_WB.instance_to_wrap.a1.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 net3258
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12501__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11667__B2 team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1653 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net3269
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\] net942
+ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and3_1
XANTENNA__08532__A1 _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08918__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18057__1433 vssd1 vssd1 vccd1 vccd1 _18057__1433/HI net1433 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ net511 _07039_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _06211_ _06141_ net504 vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08835__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ net2545 net284 net407 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
X_13490_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _05010_ vssd1 vssd1
+ vccd1 vccd1 _03843_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12441_ net2709 net200 net415 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XANTENNA__08653__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13041__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10257__A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09796__B1 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15160_ net1254 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
X_12372_ net2977 net237 net423 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08950__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14111_ net787 _04236_ _04237_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__and3_4
X_11323_ _06840_ _07586_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10945__A3 _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13568__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15091_ net1189 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04210_ _04211_ vssd1
+ vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__o21a_1
XANTENNA__13344__B2 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11254_ _06992_ _07107_ _07098_ net546 vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_28_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10205_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[1\] net737 net716 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11185_ _06211_ _06277_ _06347_ _06414_ net505 net517 vssd1 vssd1 vccd1 vccd1 _07449_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17918__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17801_ clknet_leaf_59_wb_clk_i _03358_ _01622_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_10136_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[2\] net750 _04661_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a22o_1
XANTENNA__09781__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15993_ net1355 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__inv_2
XANTENNA__11107__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13647__A2 _07510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14399__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ clknet_leaf_97_wb_clk_i _03290_ _01553_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10067_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\] net730 _06321_ _06324_
+ _06326_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a2111o_1
X_14944_ net1274 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XANTENNA__12411__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11658__B2 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18146__1520 vssd1 vssd1 vccd1 vccd1 _18146__1520/HI net1520 sky130_fd_sc_hd__conb_1
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11122__A3 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__B team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17663_ clknet_leaf_2_wb_clk_i _03223_ _01526_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14875_ net1315 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16614_ clknet_leaf_87_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[0\]
+ _00477_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13826_ team_01_WB.instance_to_wrap.cpu.c0.count\[14\] team_01_WB.instance_to_wrap.cpu.c0.count\[13\]
+ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17594_ clknet_leaf_33_wb_clk_i _03154_ _01457_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14072__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16545_ clknet_leaf_64_wb_clk_i _02173_ _00408_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _07714_ vssd1 vssd1 vccd1 vccd1
+ _04068_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10969_ _07231_ _07232_ net528 vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__mux2_1
XANTENNA__08826__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12708_ net2063 net285 net385 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16476_ clknet_leaf_109_wb_clk_i net1957 _00339_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11830__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ team_01_WB.instance_to_wrap.a1.curr_state\[0\] _04010_ vssd1 vssd1 vccd1
+ vccd1 _04011_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18215_ net1586 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15427_ net1219 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XANTENNA__13032__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ net2780 net199 net391 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XANTENNA__10167__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18146_ net1520 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
XANTENNA__09787__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16322__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15358_ net1291 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17448__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09251__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18102__1476 vssd1 vssd1 vccd1 vccd1 _18102__1476/HI net1476 sky130_fd_sc_hd__conb_1
XFILLER_0_130_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold205 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\] vssd1 vssd1 vccd1 vccd1
+ net1821 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ net1974 _04449_ net1172 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13478__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18077_ net1451 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
Xhold216 team_01_WB.instance_to_wrap.a1.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 net1832
+ sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ net1190 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold227 _02007_ vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _01983_ vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold249 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ clknet_leaf_129_wb_clk_i _02588_ _00891_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09003__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09394__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15693__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16472__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ net988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[6\] net949 vssd1
+ vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and3_1
Xfanout707 net710 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_2
Xfanout718 _04674_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 net730 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _05063_ _05064_ net578 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__mux2_2
XANTENNA__13099__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\] net915 vssd1
+ vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__and3_1
XANTENNA__13925__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11726__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12321__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[23\] net662 net624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a22o_1
XANTENNA__10630__A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11649__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08663_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\] net739 net729 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\]
+ _04916_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08594_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] net958
+ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1082_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13810__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11461__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _08022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09569__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09215_ _05468_ _05469_ _05470_ _05471_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15868__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12991__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout605_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13574__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09146_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] net617 _05381_ _05402_
+ net672 vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10388__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09077_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[18\] net642 _05311_
+ _05319_ net670 vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10805__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16815__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13326__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold750 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11337__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout974_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _02137_ vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\] vssd1 vssd1 vccd1 vccd1
+ net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 team_01_WB.instance_to_wrap.cpu.f0.num\[16\] vssd1 vssd1 vccd1 vccd1 net2410
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10243__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09979_ _06232_ _06233_ _06234_ _06235_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__or4_1
XANTENNA__13629__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12990_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[28\] net241 net361 vssd1
+ vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
Xhold1450 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3066 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08648__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1461 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net3088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11941_ net2745 net288 net471 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__mux2_1
Xhold1483 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1494 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14660_ net1373 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
X_11872_ net678 _07414_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13611_ _03815_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10823_ _05241_ _05309_ _05378_ _05448_ net503 net518 vssd1 vssd1 vccd1 vccd1 _07087_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13262__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14591_ net1371 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
X_16330_ clknet_leaf_63_wb_clk_i net1726 _00198_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10076__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13542_ net185 _07890_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _06880_ _07017_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__nor2_1
XANTENNA__09481__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08383__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ clknet_leaf_58_wb_clk_i _01898_ _00129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10685_ _06856_ _06867_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__nand2_1
X_13473_ _03813_ _03821_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a21oi_1
X_18000_ clknet_leaf_62_wb_clk_i _03549_ _01820_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15212_ net1264 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_12424_ net1887 net245 net421 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09776__A _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16192_ clknet_leaf_88_wb_clk_i _01859_ _00060_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10379__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16495__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15143_ net1195 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12406__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08441__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net2570 net302 net491 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17740__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11306_ _06664_ net334 vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__nand2_1
X_15074_ net1311 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
X_12286_ net2008 net272 net431 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux2_1
X_18044__1606 vssd1 vssd1 vccd1 vccd1 net1606 _18044__1606/LO sky130_fd_sc_hd__conb_1
XFILLER_0_103_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14025_ net1172 _04153_ _04195_ _04200_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__and4_2
XFILLER_0_43_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11237_ _06030_ _07198_ net325 vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a21o_1
XANTENNA__11879__A1 _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12930__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ _06525_ _06593_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09942__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17890__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14278__C1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ net579 _06381_ _06349_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12141__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ net1387 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__inv_2
X_11099_ _07106_ _07362_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17715_ clknet_leaf_110_wb_clk_i _03275_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09016__A _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ net1248 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11980__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17120__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17646_ clknet_leaf_55_wb_clk_i _03206_ _01509_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14858_ net1341 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XANTENNA__10854__A2 _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13809_ net486 team_01_WB.instance_to_wrap.cpu.f0.next_write_i _04478_ vssd1 vssd1
+ vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17577_ clknet_leaf_49_wb_clk_i _03137_ _01440_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14789_ net1331 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16528_ clknet_leaf_61_wb_clk_i _02156_ _00391_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17270__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__B _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16459_ clknet_leaf_100_wb_clk_i _02087_ _00322_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09000_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[19\] net609 _05247_
+ _05248_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_89_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16838__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13556__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11567__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18129_ net1503 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12316__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13308__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18056__1432 vssd1 vssd1 vccd1 vccd1 _18056__1432/HI net1432 sky130_fd_sc_hd__conb_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09902_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] net621 _06146_ _06150_
+ _06155_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 net506 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 net519 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10063__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
X_09833_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[7\] _04765_ _06072_
+ _06073_ _06093_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__a2111o_1
Xfanout548 _05651_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09852__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12051__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _05993_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nor2_1
XANTENNA__10360__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08715_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\] net691 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[23\]
+ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09695_ net582 _05958_ _05924_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a21o_1
XANTENNA__11890__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1297_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ net1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\] net931
+ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08577_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\] net648 net622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout722_A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08671__B1 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10238__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10470_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] net958
+ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ net1098 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] net862
+ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12226__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ net2589 net234 net447 vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11109__A2_N net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10781__A1 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ net2628 net239 net455 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold580 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _07285_ net322 _07158_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15830_ net1304 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__inv_2
XANTENNA__17143__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14275__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11089__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15761_ net1200 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XANTENNA__12286__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ net1026 _07478_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1280 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09151__A1 _05414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17500_ clknet_leaf_16_wb_clk_i _03060_ _01363_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14712_ net1396 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
Xhold1291 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
X_18101__1475 vssd1 vssd1 vccd1 vccd1 _18101__1475/HI net1475 sky130_fd_sc_hd__conb_1
X_11924_ net2029 net315 net476 vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
X_15692_ net1263 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17293__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ clknet_leaf_10_wb_clk_i _02991_ _01294_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13235__A0 _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ net1347 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
X_11855_ _07972_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__inv_2
XANTENNA_output105_A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__B1 _06310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13786__A1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17362_ clknet_leaf_38_wb_clk_i _02922_ _01225_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10806_ _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__inv_2
X_14574_ net1339 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11257__C_N _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11786_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] _07858_ vssd1 vssd1
+ vccd1 vccd1 _07916_ sky130_fd_sc_hd__nor2_1
XANTENNA__09454__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16313_ clknet_leaf_112_wb_clk_i _01947_ _00181_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13525_ _03755_ _03756_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__and2_1
X_10737_ net545 _06996_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__nor2_1
X_17293_ clknet_leaf_19_wb_clk_i _02853_ _01156_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13538__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16244_ clknet_leaf_79_wb_clk_i _00024_ _00112_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13456_ _03807_ _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__nand2_1
XANTENNA__09206__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10668_ _04988_ _05012_ _06872_ _06928_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__a221o_1
XANTENNA__09937__C net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08841__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ net2771 net288 net419 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16175_ clknet_leaf_90_wb_clk_i _01843_ _00043_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12136__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13387_ net2584 net327 net351 team_01_WB.instance_to_wrap.cpu.f0.i\[11\] vssd1 vssd1
+ vccd1 vccd1 _01896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10599_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _06851_ _06854_ vssd1 vssd1
+ vccd1 vccd1 _06863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XANTENNA__10221__B1 _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_15126_ net1305 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
X_12338_ net3148 net235 net490 vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11975__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15057_ net1195 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_12269_ net2884 net207 net433 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__mux2_1
XANTENNA__13710__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14008_ _04163_ _04171_ _04181_ _04188_ _04170_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a32o_1
XANTENNA__09672__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11707__C team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14266__A2 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16510__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17636__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ net1330 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__inv_2
X_08500_ net1002 net864 vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09480_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] net662 _05722_
+ _05726_ _05734_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08431_ net1131 net919 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__and2_1
XANTENNA__11723__B team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17629_ clknet_leaf_14_wb_clk_i _03189_ _01492_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16660__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _04621_ _04624_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09445__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11252__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ net3165 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[55\] net1044 vssd1 vssd1
+ vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10058__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10460__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09847__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10355__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12046__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A _07970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1045_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__B1 _04685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10763__A1 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17166__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _07984_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
Xfanout312 _07994_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
Xfanout323 net325 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_121_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout334 net336 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout672_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _06870_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08479__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_2
X_09816_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[7\] net870 vssd1
+ vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout367 net370 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_6
Xfanout378 _03570_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 _03567_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_8
XFILLER_0_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10521__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09747_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[10\] net907
+ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout937_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13605__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] net908
+ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and3_1
XANTENNA__08495__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13217__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08629_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[29\] net653 net636 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a22o_1
XANTENNA__08892__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18043__1605 vssd1 vssd1 vccd1 vccd1 net1605 _18043__1605/LO sky130_fd_sc_hd__conb_1
X_11640_ net2010 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] net840 vssd1 vssd1
+ vccd1 vccd1 _03321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11571_ _07795_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__A2 _07140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ net1859 net808 net803 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1
+ vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10522_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\] net943
+ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14290_ net1367 _04439_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13241_ _03725_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\] net829 vssd1 vssd1
+ vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
X_10453_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[26\] net763 net590 vssd1 vssd1
+ vccd1 vccd1 _06717_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input66_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[27\] net632 net611 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[27\]
+ _06644_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__a221o_1
X_13172_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[62\] net2869 net820 vssd1 vssd1
+ vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12123_ net3174 net264 net453 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
X_17980_ clknet_leaf_59_wb_clk_i _03529_ _01800_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.write_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16931_ clknet_leaf_120_wb_clk_i _02491_ _00794_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12054_ net2931 net273 net459 vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__mux2_1
XANTENNA__17659__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08389__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _07034_ _07038_ net512 vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__mux2_1
X_16862_ clknet_leaf_3_wb_clk_i _02422_ _00725_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14248__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15813_ net1225 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__inv_2
X_16793_ clknet_leaf_17_wb_clk_i _02353_ _00656_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15744_ net1286 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12956_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] net1055 net365 _03643_
+ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18055__1431 vssd1 vssd1 vccd1 vccd1 _18055__1431/HI net1431 sky130_fd_sc_hd__conb_1
XANTENNA__08836__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ net2781 net232 net477 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__mux2_1
X_15675_ net1299 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12887_ net1025 _07585_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nand2_1
XANTENNA__13759__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17414_ clknet_leaf_141_wb_clk_i _02974_ _01277_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14626_ net1410 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XANTENNA__17039__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ _07853_ _07958_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17345_ clknet_leaf_136_wb_clk_i _02905_ _01208_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14557_ net1407 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
X_11769_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] _07860_ vssd1 vssd1
+ vccd1 vccd1 _07902_ sky130_fd_sc_hd__nor2_1
XANTENNA__16127__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _03761_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17276_ clknet_leaf_14_wb_clk_i _02836_ _01139_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09667__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14488_ net1385 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10993__B2 _07185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16227_ clknet_leaf_38_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[8\]
+ _00095_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13439_ _03774_ _03791_ _03773_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a21o_1
XANTENNA__10175__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09964__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16158_ clknet_leaf_79_wb_clk_i _01826_ net1172 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10745__A1 _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15109_ net1222 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
X_08980_ net1142 net576 net577 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a21o_1
X_16089_ net1372 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__inv_2
XANTENNA__13695__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11170__A1 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14239__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ net1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\] net856 vssd1
+ vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09115__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09532_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[9\] net868 vssd1
+ vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\] net847 vssd1
+ vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout253_A _07934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08414_ net985 _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09394_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[13\] net907
+ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__and3_1
XANTENNA__09418__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08345_ net1631 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08626__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout420_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10433__B1 _06695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[80\] net2546 net1045 vssd1 vssd1
+ vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10984__A1 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15876__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10516__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16556__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18100__1474 vssd1 vssd1 vccd1 vccd1 _18100__1474/HI net1474 sky130_fd_sc_hd__conb_1
XANTENNA__10736__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17801__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_A _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12504__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11628__B _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1107 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1 vccd1
+ net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1123 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_2
Xfanout1129 net1134 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_2
XANTENNA__08157__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09354__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout186 net189 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
Xfanout197 _07869_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12810_ net1893 net252 net373 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
X_13790_ net563 _07776_ _04093_ net786 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ net1818 net284 net380 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ net1271 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
X_12672_ net3126 net198 net387 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08953__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09409__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14411_ net1308 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11623_ net497 _07826_ net2069 net839 vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__o2bb2a_1
X_15391_ net1296 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17331__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17130_ clknet_leaf_48_wb_clk_i _02690_ _00993_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10424__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14342_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1
+ vccd1 _02256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11554_ team_01_WB.instance_to_wrap.cpu.f0.i\[8\] _07739_ vssd1 vssd1 vccd1 vccd1
+ _07785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire554 _06589_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_1
X_10505_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[25\] net664 _06768_
+ net672 vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__a211o_1
X_17061_ clknet_leaf_131_wb_clk_i _02621_ _00924_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14273_ _04421_ _04423_ _04425_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__or4_1
X_11485_ net483 _07728_ net320 vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16012_ net1406 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13224_ net2279 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\] net827 vssd1 vssd1
+ vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09042__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\] net662 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__a22o_1
XANTENNA__17481__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ net2685 net2575 net824 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
X_10367_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\] net744 net698 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12414__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12106_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\] net204 net452 vssd1
+ vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__mux2_1
X_10298_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\] net963 vssd1
+ vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__and3_1
X_13086_ _05958_ _07806_ _03704_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__a21bo_1
X_17963_ clknet_leaf_85_wb_clk_i net1684 _01783_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08148__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16914_ clknet_leaf_31_wb_clk_i _02474_ _00777_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12037_ net2804 net206 net460 vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17894_ clknet_leaf_99_wb_clk_i _03444_ _01714_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[53\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10161__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16845_ clknet_leaf_16_wb_clk_i _02405_ _00708_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11554__A team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15026__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16776_ clknet_leaf_45_wb_clk_i _02336_ _00639_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _03556_ _04169_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__and2_1
XANTENNA__09648__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09024__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ net1247 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
X_12939_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] net1053 net364 _03631_
+ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16429__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15658_ net1202 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XANTENNA__09959__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14609_ net1404 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15589_ net1222 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
XANTENNA__13601__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08130_ net486 net564 net784 vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__o21a_1
X_17328_ clknet_leaf_25_wb_clk_i _02888_ _01191_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08084__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09397__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ team_01_WB.instance_to_wrap.cpu.f0.num\[22\] vssd1 vssd1 vccd1 vccd1 _04492_
+ sky130_fd_sc_hd__inv_2
XANTENNA__17824__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17259_ clknet_leaf_46_wb_clk_i _02819_ _01122_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13928__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12324__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18042__1604 vssd1 vssd1 vccd1 vccd1 net1604 _18042__1604/LO sky130_fd_sc_hd__conb_1
XFILLER_0_80_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08963_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[19\] net729 _05214_
+ _05219_ _05222_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_110_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ _05154_ _05155_ _05156_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__or4_1
XANTENNA__11143__A1 _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09860__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__A1 _07153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10779__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09515_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] net741 net702 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[9\]
+ _05774_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12994__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A _04761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09446_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\] net745 net725 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09377_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[13\] net725 net700 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08328_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[28\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[20\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ net2801 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[89\] net1048 vssd1 vssd1
+ vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
XANTENNA__11003__A1_N net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11270_ net324 _07201_ _07524_ _07533_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__o31a_1
XFILLER_0_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] net760 _06483_ _06484_
+ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__a22o_4
XFILLER_0_28_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12234__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__B2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ net581 _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__or2_1
X_10083_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] net760 _06345_ _06346_
+ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__a22o_4
X_14960_ net1256 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
Xhold9 team_01_WB.instance_to_wrap.cpu.RU0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1625
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ net2582 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[24\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14891_ net1219 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12882__B2 _03590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ clknet_leaf_105_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[16\]
+ _00493_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13842_ team_01_WB.instance_to_wrap.cpu.c0.count\[2\] team_01_WB.instance_to_wrap.cpu.c0.count\[1\]
+ team_01_WB.instance_to_wrap.cpu.c0.count\[0\] team_01_WB.instance_to_wrap.cpu.c0.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16561_ clknet_leaf_9_wb_clk_i _02189_ _00424_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13773_ net1677 net784 _04079_ _04080_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ _07161_ _07248_ net522 vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15512_ net1255 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
X_12724_ net2492 net311 net386 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XANTENNA__09779__A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16492_ clknet_leaf_108_wb_clk_i _02120_ _00355_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16721__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18231_ net1590 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ net1186 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12655_ net2136 net244 net393 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12409__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18162_ net1536 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
XANTENNA__12937__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11606_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[23\] net572 vssd1 vssd1 vccd1
+ vccd1 _07818_ sky130_fd_sc_hd__nand2_1
X_15374_ net1233 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ net2374 net263 net400 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09802__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ clknet_leaf_125_wb_clk_i _02673_ _00976_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14325_ net1703 _04459_ _04460_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__o21a_1
X_18093_ net1467 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11537_ _04476_ _07771_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16871__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10156__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1 vccd1
+ net2025 sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ clknet_leaf_7_wb_clk_i _02604_ _00907_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14256_ _04398_ _04400_ _04402_ _04411_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__or4_2
X_11468_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] net1062 _07720_ vssd1 vssd1 vccd1
+ vccd1 _07721_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ net2431 net2149 net830 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10419_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[26\] net725 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\]
+ _06669_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__a221o_1
X_14187_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\] _04263_ _04269_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__a22o_1
XANTENNA__12144__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10176__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__A1 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _04632_ _07662_ _04631_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09019__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ net2571 net2528 net820 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09318__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11983__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ net355 _03698_ _03699_ net836 net1628 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a32o_1
X_17946_ clknet_leaf_79_wb_clk_i _03496_ _01766_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16140__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1109 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11125__A1 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09869__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08526__C1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09680__C net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12873__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17877_ clknet_leaf_104_wb_clk_i _03427_ _01697_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[36\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16251__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16828_ clknet_leaf_15_wb_clk_i _02388_ _00691_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12625__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16759_ clknet_leaf_10_wb_clk_i _02319_ _00622_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09300_ net977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\] net962 vssd1
+ vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08593__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13930__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09231_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] net950
+ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12319__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09162_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[16\] net917 vssd1
+ vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08113_ team_01_WB.instance_to_wrap.cpu.f0.i\[11\] _04496_ _04500_ team_01_WB.instance_to_wrap.cpu.f0.i\[2\]
+ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09093_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[17\] net914 vssd1
+ vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10066__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_A _07943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08044_ team_01_WB.instance_to_wrap.cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1 _04475_
+ sky130_fd_sc_hd__inv_2
XANTENNA__08532__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09855__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold921 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09557__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold943 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13353__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12054__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold954 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold965 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1125_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold976 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09995_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\] net918 vssd1
+ vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__and3_1
XANTENNA__12989__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout585_A _04157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13105__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _05136_ _05203_ _05204_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__o21bai_2
Xhold1610 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1
+ net3226 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1621 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3237 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net3248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ net1128 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[21\] net954
+ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1643 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[0\] vssd1 vssd1 vccd1 vccd1
+ net3259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10810__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1654 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net3270
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10770_ _06347_ _06277_ net507 vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[12\] net748 net695 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12229__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12919__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ net3232 net286 net415 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XANTENNA__09245__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12371_ net3082 net205 net425 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ net790 net788 _04243_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__and3_4
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11322_ _04959_ _06838_ _04957_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13568__B _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15090_ net1180 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[7\] _04210_ net565 vssd1
+ vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a21boi_1
XANTENNA__13344__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11253_ _06971_ _07312_ _07320_ _06955_ _07516_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11355__B2 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[1\] net928 vssd1
+ vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__and3_1
X_11184_ _06884_ net325 _07444_ _07447_ _07443_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__o311a_1
XFILLER_0_105_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17800_ clknet_leaf_68_wb_clk_i _03357_ _01621_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.i\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_10135_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[2\] net946 vssd1
+ vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__and3_1
XANTENNA__08771__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15992_ net1381 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14943_ net1298 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
X_10066_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[3\] net952 vssd1
+ vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17731_ clknet_leaf_96_wb_clk_i _03289_ _01552_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11816__B _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08397__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14874_ net1346 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
X_17662_ clknet_leaf_13_wb_clk_i _03222_ _01525_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13825_ team_01_WB.instance_to_wrap.cpu.c0.count\[12\] _04117_ vssd1 vssd1 vccd1
+ vccd1 _04118_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16613_ clknet_leaf_86_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_read_i _00476_
+ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.READ_I sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17593_ clknet_leaf_125_wb_clk_i _03153_ _01456_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11832__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16544_ clknet_leaf_62_wb_clk_i _02172_ _00407_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ net1650 _04067_ net783 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
X_10968_ _07088_ _07093_ net509 vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__mux2_1
XANTENNA__09484__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09302__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ net2790 net222 net385 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__mux2_1
XANTENNA__08844__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18041__1603 vssd1 vssd1 vccd1 vccd1 net1603 _18041__1603/LO sky130_fd_sc_hd__conb_1
X_16475_ clknet_leaf_100_wb_clk_i _02103_ _00338_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_13687_ team_01_WB.instance_to_wrap.a1.WRITE_I team_01_WB.instance_to_wrap.a1.READ_I
+ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12139__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10899_ _06697_ _06752_ net499 vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18214_ net602 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15426_ net1292 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
X_12638_ net3150 net288 net391 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XANTENNA__09236__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11978__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18145_ net1519 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
X_15357_ net1284 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12569_ net2142 net203 net401 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] _04449_ vssd1 vssd1 vccd1
+ vccd1 _04450_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18076_ net1450 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
Xhold206 _03512_ vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ net1256 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold217 _01986_ vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold228 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17027_ clknet_leaf_119_wb_clk_i _02587_ _00890_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold239 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13335__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14239_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[14\] _04267_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\]
+ _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_2
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11897__A2 _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout719 _04672_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_6
XFILLER_0_123_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11429__D team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ net1110 net763 net590 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a21o_1
XANTENNA__13494__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12602__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _06031_ _06041_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__or3_1
XANTENNA__13099__B2 _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08588__A _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\] net646 net637 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[23\]
+ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17929_ clknet_leaf_101_wb_clk_i _03479_ _01749_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10630__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08514__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 net1292 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08662_ _04922_ _04923_ _04924_ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__or4_1
XANTENNA__10321__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08593_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\] net942 vssd1
+ vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11461__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12049__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10358__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1075_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\] net643 _05477_
+ net671 vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13940__A_N net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14220__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13669__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ _05405_ _05406_ _05407_ _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__or4_2
XFILLER_0_60_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1242_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10388__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09076_ _05336_ _05337_ _05338_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__or4_2
XANTENNA__08450__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13326__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold740 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10524__C net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold762 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold773 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__D1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 net2400
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 team_01_WB.instance_to_wrap.cpu.c0.count\[6\] vssd1 vssd1 vccd1 vccd1 net2411
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_89_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12512__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[5\] net639 _06241_ net672
+ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08498__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10560__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[21\] _04759_ _05174_
+ _05178_ _05180_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11636__B _07806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1440 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1451 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3067 sky130_fd_sc_hd__dlygate4sd3_1
X_11940_ net1979 net230 net471 vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1462 team_01_WB.instance_to_wrap.cpu.f0.state\[2\] vssd1 vssd1 vccd1 vccd1 net3078
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10312__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1473 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[41\] vssd1 vssd1 vccd1 vccd1
+ net3089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1484 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1495 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\] vssd1 vssd1 vccd1 vccd1
+ net3111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11871_ _07849_ _07985_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__or2_1
XANTENNA__10967__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13610_ _03822_ _03946_ _03818_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__o21a_1
X_10822_ _05241_ _05309_ net502 vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__mux2_1
X_14590_ net1409 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _03763_ _03859_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ _06485_ net505 vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11812__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16260_ clknet_leaf_71_wb_clk_i _01897_ _00128_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.num\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13472_ _03816_ _03818_ _03822_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a31o_1
XANTENNA__17072__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ _04851_ _04828_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__nand2b_1
XANTENNA__14211__B1 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15211_ net1204 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XANTENNA__13579__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ net2489 net316 net419 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__mux2_1
X_16191_ clknet_leaf_88_wb_clk_i _01858_ _00059_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10379__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15142_ net1287 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12354_ net2598 net262 net491 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13317__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _06722_ _07128_ _06940_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15073_ net1312 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12285_ net2003 net246 net431 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__mux2_1
X_14024_ _04195_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nand2_2
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ _06030_ _07198_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__nor2_1
XANTENNA__12930__B _07223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13518__S net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ _06525_ _06880_ net325 vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12422__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10551__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ net579 _06381_ _06349_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__o21a_2
XANTENNA__08839__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ net1335 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__inv_2
X_11098_ _07208_ _07361_ net534 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17714_ clknet_leaf_110_wb_clk_i _03274_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10049_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\] net667 _06310_ _06312_
+ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__o22a_4
X_14926_ net1228 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17645_ clknet_leaf_50_wb_clk_i _03205_ _01508_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14857_ net1354 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ net1675 _04107_ net783 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14788_ net1331 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
X_17576_ clknet_leaf_62_wb_clk_i _03136_ _01439_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08347__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16527_ clknet_leaf_59_wb_clk_i _02155_ _00390_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13739_ net563 _04053_ _04054_ net485 vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09967__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16458_ clknet_leaf_107_wb_clk_i net2870 _00321_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14202__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13556__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13489__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15409_ net1195 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
X_16389_ clknet_leaf_70_wb_clk_i _02017_ _00252_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17565__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18128_ net1502 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
XFILLER_0_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13308__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18059_ net1435 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_09901_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[6\] net615 _06145_ _06147_
+ _06159_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_111_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout505 net506 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout516 net519 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_4
X_09832_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\] net625 _06076_ _06081_
+ _06082_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08735__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_2
Xfanout538 net540 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XANTENNA__10641__A _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14269__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _04714_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09763_ net581 net557 _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout283_A _07920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[23\] net738 net689 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09694_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] net667 _05952_ _05957_
+ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__o22a_2
XFILLER_0_59_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08645_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[28\] net954
+ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout450_A _08019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1192_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11472__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08576_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] net640 net631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_136_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10519__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08671__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13399__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12507__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11558__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09128_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] net849
+ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16932__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[18\] net851
+ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12070_ net2046 net206 net457 vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
Xhold570 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[122\] vssd1 vssd1 vccd1 vccd1
+ net2208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11021_ _05138_ _07157_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__nor2_1
XANTENNA__08726__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09117__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15760_ net1253 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
X_12972_ net1637 net606 net588 _03655_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a22o_1
XANTENNA__08956__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 team_01_WB.instance_to_wrap.a1.ADR_I\[29\] vssd1 vssd1 vccd1 vccd1 net2886
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ net1408 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
Xhold1281 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ net1944 net303 net476 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
Xhold1292 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ net1207 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__10697__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14642_ net1409 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
X_17430_ clknet_leaf_32_wb_clk_i _02990_ _01293_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13235__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11854_ _07851_ _07971_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10805_ net549 net525 vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17361_ clknet_leaf_24_wb_clk_i _02921_ _01224_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14573_ net1366 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11785_ net1977 net222 net481 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__mux2_1
XANTENNA__17588__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16312_ clknet_leaf_111_wb_clk_i _01946_ _00180_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13524_ net967 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[30\] _03874_ _03875_
+ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a22o_1
X_17292_ clknet_leaf_45_wb_clk_i _02852_ _01155_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10736_ net542 _06967_ _06997_ _06994_ _06977_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a311o_1
XFILLER_0_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16243_ clknet_leaf_79_wb_clk_i _00023_ _00111_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_13455_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _05853_ vssd1 vssd1 vccd1
+ vccd1 _03808_ sky130_fd_sc_hd__or2_1
XANTENNA__12417__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ _06877_ _06930_ _05015_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ net3168 net231 net421 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16174_ clknet_leaf_58_wb_clk_i _01842_ _00042_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13386_ net2325 net328 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1
+ vccd1 vccd1 _01897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[1\] _06851_ _06854_ vssd1 vssd1
+ vccd1 vccd1 _06862_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10221__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ net1174 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XANTENNA__08965__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_105_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12337_ net2960 net205 net492 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_121_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12941__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15056_ net1247 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12268_ net2941 net190 net431 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__mux2_1
XANTENNA__09953__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ _04170_ _04188_ _04190_ _04167_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
XANTENNA__08717__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ _06041_ _06899_ _06912_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12152__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net2833 net211 net446 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XANTENNA__09027__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11991__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15958_ net1321 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09142__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ net1281 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08350__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15889_ net1353 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16805__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ net1141 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\] net914
+ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__and3_1
XANTENNA__10400__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17628_ clknet_leaf_14_wb_clk_i _03188_ _01491_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11237__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13777__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _04621_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17559_ clknet_leaf_10_wb_clk_i _03119_ _01422_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12985__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09697__A _05923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08292_ net2401 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[56\] net1039 vssd1 vssd1
+ vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16955__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12327__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1038_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 _07970_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08708__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12062__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 _07994_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10515__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_4
Xfanout346 _06869_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_4
Xfanout357 _03670_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_4
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[7\] net870 vssd1
+ vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and3_1
Xfanout368 net370 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_6
XANTENNA__12997__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout379 net382 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_6
XANTENNA_fanout665_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[10\] net896
+ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09677_ net1016 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\] net869
+ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout832_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08495__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\] net643 net617 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[29\]
+ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17730__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\] net725 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__a22o_1
XANTENNA__11779__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12976__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13621__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ _04482_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10521_ net971 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\] net935 vssd1
+ vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09400__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12237__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11141__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13240_ _03724_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\] net831 vssd1 vssd1
+ vccd1 vccd1 _02018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] net666 _06706_ _06715_
+ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__o22a_4
XFILLER_0_33_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[63\] net2715 net825 vssd1 vssd1
+ vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
X_10383_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\] net659 _04745_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12122_ net1987 net268 net454 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__mux2_1
XANTENNA_input59_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ net2815 net248 net461 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__mux2_1
X_16930_ clknet_leaf_0_wb_clk_i _02490_ _00793_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10506__A2 _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _05138_ net340 net339 _05136_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12900__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09372__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ clknet_leaf_14_wb_clk_i _02421_ _00724_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout880 _04746_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08580__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15812_ net1269 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__inv_2
Xfanout891 net895 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12700__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ clknet_leaf_25_wb_clk_i _02352_ _00655_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15743_ net1298 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
X_12955_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[8\] _07379_ net1033 vssd1 vssd1
+ vccd1 vccd1 _03643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ net3173 net234 net475 vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12886_ net1773 net607 net589 _03593_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a22o_1
X_15674_ net1259 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16978__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17413_ clknet_leaf_132_wb_clk_i _02973_ _01276_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14625_ net1401 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
X_11837_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] _07852_ vssd1 vssd1
+ vccd1 vccd1 _07958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10159__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14556_ net1335 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17344_ clknet_leaf_141_wb_clk_i _02904_ _01207_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11768_ net2339 net288 net479 vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ _03766_ _03767_ _03856_ _03765_ _03763_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a311o_1
XANTENNA__16208__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _06978_ _06981_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__or2_2
X_17275_ clknet_leaf_36_wb_clk_i _02835_ _01138_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12147__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14487_ net1358 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ _04719_ _05243_ _06850_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__or3_2
XFILLER_0_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16226_ clknet_leaf_38_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[7\]
+ _00094_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_13438_ _03777_ _03790_ _03776_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11986__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13767__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ net1383 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__inv_2
XANTENNA__08938__A2 _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ net2451 net329 net353 team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1
+ vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ net1226 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16088_ net1376 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__inv_2
XANTENNA__09683__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15039_ net1294 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XANTENNA__13695__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08571__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\] net860 vssd1
+ vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12610__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13933__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] net882 vssd1
+ vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\] net868
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__and3_1
X_08413_ net1148 net1150 net1152 net1154 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__nor4_2
XFILLER_0_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09393_ net995 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] net871 vssd1
+ vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08344_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[4\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09858__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10433__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09220__A _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ net3094 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[73\] net1049 vssd1 vssd1
+ vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
XANTENNA__12057__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17133__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout413_A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1155_A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10984__A2 _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__A2 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__B _06348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A2 _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09593__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout782_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1108 net1110 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_2
XANTENNA__13686__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1119 net1123 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_2
XANTENNA__09890__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09354__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12520__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout198 net199 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] net760 _05991_ _05992_
+ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ net2385 net222 net380 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11863__A1_N net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ net2705 net288 net387 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14410_ net1340 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11622_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[15\] net573 vssd1 vssd1 vccd1
+ vccd1 _07826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15390_ net1315 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14341_ net2153 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09130__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11553_ team_01_WB.instance_to_wrap.cpu.f0.i\[10\] _07745_ _07782_ _07784_ vssd1
+ vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10504_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] _04741_ net621
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\] vssd1 vssd1 vccd1 vccd1
+ _06768_ sky130_fd_sc_hd__a22o_1
XANTENNA__10707__C _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17060_ clknet_leaf_138_wb_clk_i _02620_ _00923_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14166__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14272_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[111\] _04256_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[95\]
+ _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__a221o_1
Xwire555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_1
X_11484_ _07730_ _07735_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16500__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16011_ net1386 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13223_ net3244 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[19\] net831 vssd1 vssd1
+ vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] net652 net609 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[26\]
+ _06698_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13154_ net1956 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[88\] net817 vssd1 vssd1
+ vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[27\] net754 _06618_
+ _06620_ _06621_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12105_ net2839 net241 net451 vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
X_13085_ net354 _03709_ _03710_ net834 net2113 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a32o_1
X_17962_ clknet_leaf_80_wb_clk_i net1822 _01782_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16650__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10297_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\] net919 vssd1
+ vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09345__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16913_ clknet_leaf_23_wb_clk_i _02473_ _00776_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12036_ net2189 net193 net459 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17893_ clknet_leaf_104_wb_clk_i _03443_ _01713_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[52\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11152__A2 _06983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16844_ clknet_leaf_44_wb_clk_i _02404_ _00707_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12430__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16775_ clknet_leaf_133_wb_clk_i _02335_ _00638_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13987_ _04164_ _04173_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__nand2_1
X_15726_ net1230 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
X_12938_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[13\] _07551_ net1026 vssd1 vssd1
+ vccd1 vccd1 _03631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10663__A1 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15657_ net1228 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
X_12869_ _04510_ _03580_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor2_1
XANTENNA__17156__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15042__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ net1406 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08355__S net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__C net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15588_ net1270 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ clknet_leaf_18_wb_clk_i _02887_ _01190_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14539_ net1322 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14881__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ team_01_WB.instance_to_wrap.cpu.f0.num\[26\] vssd1 vssd1 vccd1 vccd1 _04491_
+ sky130_fd_sc_hd__inv_2
XANTENNA__14157__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17258_ clknet_leaf_48_wb_clk_i _02818_ _01121_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16209_ clknet_leaf_117_wb_clk_i _01876_ _00077_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13497__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17189_ clknet_leaf_132_wb_clk_i _02749_ _01052_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12605__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13928__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap855 _04760_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08792__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] net731 net720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10352__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11679__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\] net732 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12340__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__A2 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12340__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08757__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_A _03665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ _05771_ _05775_ _05776_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09445_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[12\] net687 _05694_
+ _05696_ _05701_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout530_A _06451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_A _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1272_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09376_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] net727 net721 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\]
+ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16523__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17649__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08327_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[29\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[21\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09885__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08258_ net1798 net2259 net1047 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout997_A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13356__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08189_ _04551_ _04581_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16673__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12515__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17799__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10220_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[1\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11382__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] net765 _04723_ net1110 vssd1
+ vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17029__CLK clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10082_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[3\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13910_ net3269 net794 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[23\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12250__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ net1201 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12882__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ net2170 _04111_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17179__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13772_ net484 _07712_ _07764_ net786 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a31o_1
X_16560_ clknet_leaf_7_wb_clk_i _02188_ _00423_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ _05099_ _05241_ _05309_ _05378_ net502 net516 vssd1 vssd1 vccd1 vccd1 _07248_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15511_ net1247 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
X_12723_ net2112 net259 net386 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16491_ clknet_leaf_101_wb_clk_i net1664 _00354_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18230_ net601 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12654_ net3221 net315 net391 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15442_ net1175 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
XANTENNA__09498__C net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ net496 _07817_ net2397 net838 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13595__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18161_ net1535 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
X_15373_ net1214 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
X_12585_ net2768 net267 net402 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17112_ clknet_leaf_28_wb_clk_i _02672_ _00975_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11536_ team_01_WB.instance_to_wrap.cpu.f0.i\[8\] net1065 vssd1 vssd1 vccd1 vccd1
+ _07771_ sky130_fd_sc_hd__nand2_1
XANTENNA__14139__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14324_ net1703 _04459_ net1362 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18092_ net1466 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_83_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17043_ clknet_leaf_51_wb_clk_i _02603_ _00906_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14255_ _04404_ _04406_ _04408_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__or4_1
X_11467_ _04467_ _07719_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__nor2_1
XANTENNA__12425__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[28\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[36\]
+ net821 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
X_10418_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\] net720 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__a22o_1
X_14186_ _04153_ _04344_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11398_ _07023_ _07654_ _07661_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13137_ net1633 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\] net828 vssd1 vssd1
+ vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10349_ _05138_ _05206_ _06610_ _05210_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__o31a_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10172__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\] net1031 vssd1 vssd1 vccd1
+ vccd1 _03699_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17945_ clknet_leaf_102_wb_clk_i _03495_ _01765_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09961__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11125__A2 _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ net1840 net276 net464 vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XANTENNA__12160__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17876_ clknet_leaf_75_wb_clk_i net3114 _01696_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12873__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16827_ clknet_leaf_37_wb_clk_i _02387_ _00690_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16758_ clknet_leaf_29_wb_clk_i _02318_ _00621_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15709_ net1280 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
X_16689_ clknet_leaf_55_wb_clk_i _02249_ _00552_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09230_ net974 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[15\] net953 vssd1
+ vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09161_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[16\] net930
+ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16696__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08112_ _04470_ team_01_WB.instance_to_wrap.cpu.f0.num\[18\] _04494_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17941__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09092_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[17\] net938 vssd1
+ vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ net1064 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold900 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12335__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold911 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout209_A _07879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold922 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold933 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold944 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold955 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[96\] vssd1 vssd1 vccd1 vccd1
+ net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 net2582
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold977 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09994_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] net946 vssd1
+ vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold988 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1118_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09309__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13674__B _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _05013_ _05068_ _05014_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout480_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1600 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3216 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08517__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1611 _04145_ vssd1 vssd1 vccd1 vccd1 net3227 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17321__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3238 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ net1126 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\] net931
+ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1633 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[4\] vssd1 vssd1 vccd1 vccd1
+ net3260 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08098__A2_N team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1655 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 net3271
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout745_A _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08784__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13813__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17471__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09428_ net1122 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\] net929
+ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[13\] net926 vssd1
+ vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12370_ net2901 net240 net425 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
XANTENNA__09796__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08950__C net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11321_ net322 _07583_ _07584_ net344 _07581_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__o221a_2
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12245__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _04210_ net566 _04209_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__and3b_1
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11252_ _05486_ net343 _07514_ _07515_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10203_ net1139 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[1\] net955 vssd1
+ vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__and3_1
XANTENNA__08756__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__A2 _07019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11183_ _06972_ _07139_ _07446_ _06454_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08959__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[2\] net923 vssd1
+ vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15991_ net1327 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__inv_2
XANTENNA__09781__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12304__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17730_ clknet_leaf_97_wb_clk_i _03288_ _01551_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.CU0.opcode\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_10065_ net990 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[3\] net955 vssd1
+ vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__and3_1
X_14942_ net1287 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ clknet_leaf_127_wb_clk_i _03221_ _01524_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14873_ net1380 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
X_16612_ clknet_leaf_87_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_write_i
+ _00475_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.WRITE_I sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ team_01_WB.instance_to_wrap.cpu.c0.count\[10\] team_01_WB.instance_to_wrap.cpu.c0.count\[11\]
+ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13804__A1 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17592_ clknet_leaf_27_wb_clk_i _03152_ _01455_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08694__A _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16543_ clknet_leaf_64_wb_clk_i _02171_ _00406_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ _04064_ _04066_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__nand2_1
X_10967_ _07086_ _07089_ net510 vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12706_ net2622 net226 net383 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16474_ clknet_leaf_107_wb_clk_i net2719 _00337_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_13686_ net968 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _04008_ _04009_
+ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
X_10898_ _04935_ _06643_ net499 vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ net602 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15425_ net1291 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ net2657 net233 net393 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10167__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15320__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18144_ net1518 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
X_15356_ net1235 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ net2378 net238 net401 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__mux2_1
XANTENNA__09787__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11519_ _04469_ _07731_ _07757_ _07759_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__a31o_1
X_14307_ net1366 _04448_ _04449_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nor3_1
XFILLER_0_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18075_ net1449 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XANTENNA__12155__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12499_ net2175 net195 net407 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
X_15287_ net1246 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[0\] vssd1 vssd1 vccd1 vccd1
+ net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17026_ clknet_leaf_143_wb_clk_i _02586_ _00889_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold229 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] _04253_ _04279_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\]
+ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__a22o_1
XANTENNA__08747__A0 _05009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13740__B1 _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[59\] _04253_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__a22o_1
XANTENNA__17344__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10554__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13099__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15990__A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] net644 net614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ clknet_leaf_101_wb_clk_i net2762 _01748_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[87\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1280 net1285 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_4
Xfanout1291 net1292 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08661_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[28\] net704 _04911_
+ _04912_ _04915_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a2111o_1
X_17859_ clknet_leaf_80_wb_clk_i _03409_ _01679_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_08592_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\] net958 vssd1
+ vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11282__A1 _07184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09213_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[16\] net653 net630 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1068_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[17\] net657 _05385_
+ _05390_ _05393_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13669__B _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[18\] net644 _05315_
+ _05317_ _05330_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12065__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10793__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08450__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold730 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout695_A _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold763 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08202__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold774 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1402_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[64\] vssd1 vssd1 vccd1 vccd1
+ net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09977_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[5\] net651 net636 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout862_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08498__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08928_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[21\] _04767_ _05169_
+ _05181_ _05185_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a2111o_1
Xhold1430 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 net3046
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10848__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1452 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1463 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[43\] vssd1 vssd1 vccd1 vccd1
+ net3079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08859_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[20\] net637 _05100_
+ _05107_ _05109_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__a2111o_1
Xhold1474 team_01_WB.instance_to_wrap.cpu.DM0.state\[2\] vssd1 vssd1 vccd1 vccd1 net3090
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1485 team_01_WB.instance_to_wrap.cpu.f0.num\[15\] vssd1 vssd1 vccd1 vccd1 net3101
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10943__S1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] _07848_ vssd1 vssd1 vccd1
+ vccd1 _07985_ sky130_fd_sc_hd__nor2_1
Xhold1496 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net3112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10821_ net543 _07084_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__nor2_1
XANTENNA__09403__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13262__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11144__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13540_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _03888_ net1066 vssd1
+ vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
X_10752_ _06414_ _06347_ net507 vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17217__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13471_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _05550_ _03823_ vssd1
+ vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__a21o_1
X_10683_ _06943_ _06946_ _04854_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15210_ net1199 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
X_12422_ net3035 net302 net420 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16190_ clknet_leaf_91_wb_clk_i _01857_ _00058_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08977__B1 _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16241__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15141_ net1225 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
X_12353_ net2638 net266 net493 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10784__A0 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17367__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08441__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ _07563_ _07564_ _07567_ _07562_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__o211a_1
X_15072_ net1273 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12284_ net2670 net277 net432 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14023_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__inv_2
XANTENNA__13722__B1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ net345 _07497_ _07498_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__or3b_1
XANTENNA__12703__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16391__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _06525_ net343 _07256_ _06971_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10117_ _06377_ _06379_ net574 _06350_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__a31oi_4
X_15974_ net1334 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__inv_2
X_11097_ _07358_ _07360_ net529 vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10839__A1 _06989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17713_ clknet_leaf_110_wb_clk_i _03273_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_14925_ net1216 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
X_10048_ _06303_ _06304_ _06305_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__or4_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold90 net150 vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08901__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17644_ clknet_leaf_44_wb_clk_i _03204_ _01507_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14856_ net1351 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08855__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ net564 _07771_ _04106_ net485 _04477_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a32o_1
XANTENNA__13789__B1 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17575_ clknet_leaf_126_wb_clk_i _03135_ _01438_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14787_ net1333 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ net2443 net290 net468 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10067__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16526_ clknet_leaf_57_wb_clk_i _02154_ _00389_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13738_ team_01_WB.instance_to_wrap.cpu.f0.i\[23\] _07752_ vssd1 vssd1 vccd1 vccd1
+ _04054_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11989__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16457_ clknet_leaf_99_wb_clk_i _02085_ _00320_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[69\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_89_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13669_ net772 _07414_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__nand2_1
XANTENNA__08680__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15408_ net1262 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
X_16388_ clknet_leaf_75_wb_clk_i _02016_ _00251_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11567__A2 _07734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08968__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18127_ net1501 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
X_15339_ net1204 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10194__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18058_ net1434 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_83_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09900_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[6\] net636 _06144_ _06156_
+ _06160_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__a2111o_1
X_17009_ clknet_leaf_23_wb_clk_i _02569_ _00872_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12613__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10922__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13936__C team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_4
XANTENNA__09932__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] net665 _06078_ _06080_
+ _06084_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout528 _06451_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_2
XFILLER_0_67_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09762_ team_01_WB.instance_to_wrap.cpu.CU0.bit30 net591 net581 vssd1 vssd1 vccd1
+ vccd1 _06026_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10360__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ _04974_ _04975_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__or3_1
X_09693_ _05953_ _05954_ _05955_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net982 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[28\] net931 vssd1
+ vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11472__B team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[30\] net633 net618 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[30\]
+ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout443_A _08020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1185_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16264__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A _04776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09596__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09127_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[17\] net898 vssd1
+ vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_105_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10766__A0 _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\] net897 vssd1
+ vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09893__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold560 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12523__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold571 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11020_ _07267_ _07268_ _07283_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__nor3_1
Xhold582 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[62\] vssd1 vssd1 vccd1 vccd1
+ net2198 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold593 _02138_ vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11647__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12971_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] net1055 _03582_ _03654_
+ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a22o_1
Xhold1260 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ net1377 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
Xhold1271 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11494__A1 _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ net2291 net263 net476 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__mux2_1
Xhold1293 team_01_WB.instance_to_wrap.cpu.K0.code\[1\] vssd1 vssd1 vccd1 vccd1 net2909
+ sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ net1196 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14641_ net1386 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _07850_ vssd1 vssd1 vccd1
+ vccd1 _07971_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10049__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17360_ clknet_leaf_23_wb_clk_i _02920_ _01223_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _07056_ _07057_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14572_ net1340 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
X_11784_ net775 _07912_ _07913_ _07914_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_71_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16311_ clknet_leaf_111_wb_clk_i _01945_ _00179_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13523_ net767 _07082_ net1066 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o21a_1
X_17291_ clknet_leaf_46_wb_clk_i _02851_ _01154_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ _06967_ _06997_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16242_ clknet_leaf_79_wb_clk_i _00022_ _00110_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14196__B1 _04258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ _05069_ _06876_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__nand2_1
X_13454_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] _05853_ vssd1 vssd1 vccd1
+ vccd1 _03807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12405_ net3170 net235 net419 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13385_ net2218 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1
+ vccd1 vccd1 _01898_ sky130_fd_sc_hd__a22o_1
X_16173_ clknet_leaf_58_wb_clk_i _01841_ _00041_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10757__A0 _07011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10597_ _06853_ _06859_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15124_ net1243 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
X_12336_ net2752 net239 net492 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__B _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12433__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ net3051 net196 net433 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__mux2_1
X_15055_ net1251 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14214__A _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14006_ _04163_ _03556_ _04181_ _03557_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__a31o_1
XANTENNA__09375__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _05890_ _07370_ _06043_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__a21o_1
X_12198_ net2913 net291 net444 vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
X_11149_ _07397_ net324 _07345_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14120__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13930__A_N net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ net1330 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__inv_2
X_14908_ net1277 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15888_ net1353 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__inv_2
X_17627_ clknet_leaf_36_wb_clk_i _03187_ _01490_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14839_ net1339 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XANTENNA__10189__A _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08360_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[3\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[2\]
+ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[1\] team_01_WB.instance_to_wrap.cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and4b_2
X_17558_ clknet_leaf_32_wb_clk_i _03118_ _01421_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08882__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08102__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08102__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_114_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_3_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16509_ clknet_leaf_78_wb_clk_i net2388 _00372_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12985__A1 team_01_WB.instance_to_wrap.a1.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18195__1569 vssd1 vssd1 vccd1 vccd1 _18195__1569/HI net1569 sky130_fd_sc_hd__conb_1
X_08291_ net3160 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[57\] net1049 vssd1 vssd1
+ vccd1 vccd1 _03456_ sky130_fd_sc_hd__mux2_1
X_17489_ clknet_leaf_20_wb_clk_i _03049_ _01352_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12608__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14187__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10460__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12737__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10748__A0 _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10355__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10212__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11748__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12343__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09218__A _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _07970_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout314 net317 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_2
Xfanout325 _06949_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout393_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _06984_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_4
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09814_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[7\] net844 vssd1
+ vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__and3_1
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_2
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1100_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10090__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[10\] net886
+ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout658_A _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ net1095 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\] net883
+ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__and3_1
XANTENNA__08268__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[29\] net623 net611 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08892__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout825_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08558_ _04818_ _04819_ _04820_ _04821_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12976__B2 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ net1084 net864 vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__and2_4
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12518__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14178__B1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ net973 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[24\] net928 vssd1
+ vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10451_ _06708_ _06710_ _06712_ _06714_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10265__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\] net2202 net818 vssd1 vssd1
+ vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
X_10382_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[27\] _04741_ net645
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\] vssd1 vssd1 vccd1 vccd1
+ _06646_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12121_ net2742 net273 net451 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__mux2_1
XANTENNA__12253__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12052_ net2302 net275 net461 vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XANTENNA__09128__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08032__A team_01_WB.instance_to_wrap.cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11164__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ net332 _05137_ _05135_ net334 vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13873__A team_01_WB.instance_to_wrap.cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12900__B2 _03603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16860_ clknet_leaf_16_wb_clk_i _02420_ _00723_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout870 _04750_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
XANTENNA__09109__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15811_ net1221 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__inv_2
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_4
Xfanout892 net895 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_2
X_16791_ clknet_leaf_10_wb_clk_i _02351_ _00654_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_15742_ net1288 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
X_12954_ net1829 net606 net588 _03642_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
Xhold1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11905_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[27\] net204 net477 vssd1
+ vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__mux2_1
X_15673_ net1192 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
X_12885_ net366 _03591_ _03592_ net1056 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17412_ clknet_leaf_138_wb_clk_i _02972_ _01275_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14624_ net1406 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
X_11836_ net2377 net273 net479 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17343_ clknet_leaf_1_wb_clk_i _02903_ _01206_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14555_ net1408 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12428__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08635__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net774 _07900_ _07899_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__a21o_2
XANTENNA__10737__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11416__A1_N net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14169__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ _03766_ _03767_ _03856_ _03765_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a31o_1
X_17274_ clknet_leaf_36_wb_clk_i _02834_ _01137_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10718_ _06978_ _06981_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ net1358 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
X_11698_ net3143 net152 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16225_ clknet_leaf_42_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[6\]
+ _00093_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13437_ _03787_ _03788_ _03779_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__a21o_1
X_10649_ _05822_ _05788_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__and2b_1
XANTENNA__10175__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13392__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16156_ net1383 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__inv_2
X_13368_ net2425 net328 net352 team_01_WB.instance_to_wrap.cpu.f0.i\[30\] vssd1 vssd1
+ vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09964__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15107_ net1222 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12163__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net2114 net270 net427 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
X_16087_ net1366 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__inv_2
XANTENNA__10472__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299_ net125 net810 net805 net1668 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15038_ net1312 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XANTENNA__13783__A team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08877__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16989_ clknet_leaf_127_wb_clk_i _02549_ _00852_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ net998 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\] net891 vssd1
+ vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09461_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] net882
+ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__and3_1
XANTENNA__16922__CLK clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08412_ net978 net919 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__and2_4
XFILLER_0_87_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09392_ net994 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[13\] net904 vssd1
+ vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09501__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08343_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[5\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12338__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ net2058 net2019 net1052 vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10433__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10984__A3 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1050_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout406_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1148_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17428__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11478__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13686__A2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_1
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13693__A team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16452__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17578__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12801__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout942_A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout199 net201 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09728_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[10\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09511__B1 _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09659_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[11\] net760 _05921_ _05922_
+ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12670_ net2537 net230 net389 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08953__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__A1 _07510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11621_ net497 _07825_ net2315 net839 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_120_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12248__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14340_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[18\] vssd1 vssd1 vccd1
+ vccd1 _02258_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10424__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _04475_ _07704_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11621__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[25\] net616 net613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\]
+ _06766_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11483_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] net1061 _07727_ _07734_ team_01_WB.instance_to_wrap.cpu.f0.i\[30\]
+ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__a41o_1
XFILLER_0_80_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14271_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[79\] _04246_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[71\]
+ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire556 _06069_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_1
X_16010_ net1394 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__inv_2
XANTENNA__09578__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input71_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[26\] net629 net624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__a22o_1
X_13222_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[12\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[20\]
+ net823 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XANTENNA__13374__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09042__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ net2862 net2347 net828 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10365_ _06619_ _06626_ _06627_ _06628_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12104_ net2676 net207 net452 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
X_13084_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\] net1028 vssd1 vssd1 vccd1
+ vccd1 _03710_ sky130_fd_sc_hd__or2_1
XANTENNA__11137__A0 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17961_ clknet_leaf_106_wb_clk_i net1681 _01781_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_10296_ net581 _06559_ _06526_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16912_ clknet_leaf_30_wb_clk_i _02472_ _00775_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12035_ net2579 net194 net460 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
X_17892_ clknet_leaf_75_wb_clk_i _03442_ _01712_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12885__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12711__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18194__1568 vssd1 vssd1 vccd1 vccd1 _18194__1568/HI net1568 sky130_fd_sc_hd__conb_1
XANTENNA__08697__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16843_ clknet_leaf_56_wb_clk_i _02403_ _00706_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16945__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16774_ clknet_leaf_139_wb_clk_i _02334_ _00637_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13986_ _04160_ _04164_ _04172_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15725_ net1216 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
X_12937_ net1734 net605 net587 _03630_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09024__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15656_ net1183 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
X_12868_ net1034 _03578_ _03579_ net1161 vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__a211o_1
XANTENNA__09959__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14607_ net1372 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
X_11819_ net2995 net215 net479 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XANTENNA__13062__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ net1222 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XANTENNA__12158__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12799_ net2717 net240 net373 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XANTENNA__13601__A2 _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17326_ clknet_leaf_51_wb_clk_i _02886_ _01189_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14538_ net1318 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17257_ clknet_leaf_42_wb_clk_i _02817_ _01120_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14469_ net1336 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16208_ clknet_leaf_116_wb_clk_i _01875_ _00076_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17188_ clknet_leaf_129_wb_clk_i _02748_ _01051_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09033__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16139_ net1314 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09991__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08961_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[19\] net738 net705 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12876__A0 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12621__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\] net719 net706 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\]
+ _05148_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11143__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08400__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09513_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] net746 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09444_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[12\] net733 net701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[12\]
+ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09231__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13053__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09375_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[13\] net697 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout523_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1265_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08326_ net2640 net2552 net1041 vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08257_ net2482 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[91\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03490_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16818__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13356__A1 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ _04553_ _04575_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11367__A0 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout892_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13108__A1 _06450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] net760 _06412_ _06413_
+ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__a22o_2
XANTENNA__09980__B1 _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A0 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16968__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10081_ _06336_ _06337_ _06342_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__or4_2
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09406__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18069__1443 vssd1 vssd1 vccd1 vccd1 _18069__1443/HI net1443 sky130_fd_sc_hd__conb_1
X_13840_ _04114_ _04126_ _04129_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.next_count\[7\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__10893__A2 _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ _07712_ _07774_ _04014_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] net563
+ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10983_ _05419_ _06920_ _06925_ _07227_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15510_ net1258 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
X_12722_ net2576 net300 net386 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16490_ clknet_leaf_102_wb_clk_i _02118_ _00353_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11390__B _07585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15441_ net1193 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XANTENNA__13044__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ net3092 net304 net392 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18160_ net1534 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
X_11604_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[24\] net572 vssd1 vssd1 vccd1
+ vccd1 _07817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ net1252 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_142_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12584_ net2376 net272 net399 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__mux2_1
X_17111_ clknet_leaf_10_wb_clk_i _02671_ _00974_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14323_ net1362 _04458_ _04459_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nor3_1
XANTENNA__10802__C1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18091_ net1465 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_11535_ team_01_WB.instance_to_wrap.cpu.f0.i\[6\] team_01_WB.instance_to_wrap.cpu.f0.i\[5\]
+ _07769_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__and3_1
XANTENNA__16498__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12706__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17743__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09287__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17042_ clknet_leaf_31_wb_clk_i _02602_ _00905_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14254_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[126\] _04275_ _04280_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\]
+ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11466_ team_01_WB.instance_to_wrap.cpu.f0.i\[21\] _07718_ vssd1 vssd1 vccd1 vccd1
+ _07719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10734__B _06995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[29\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[37\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\] net749 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14185_ _04238_ _04273_ _04343_ _04287_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__nor4b_1
X_11397_ _07600_ _07655_ _07659_ _07660_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ net1640 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[106\] net827 vssd1 vssd1
+ vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
X_10348_ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__inv_2
XANTENNA__09019__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17893__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15318__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _06530_ _06534_ _06538_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13067_ _03666_ _03697_ net1027 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12441__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ clknet_leaf_101_wb_clk_i _03494_ _01764_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11125__A3 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12018_ net2985 net215 net463 vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XANTENNA__08858__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17875_ clknet_leaf_80_wb_clk_i _03425_ _01695_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16826_ clknet_leaf_35_wb_clk_i _02386_ _00689_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16757_ clknet_leaf_8_wb_clk_i _02317_ _00620_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13283__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\] _04158_ _04161_ net1171
+ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__o211a_1
X_15708_ net1278 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ clknet_leaf_54_wb_clk_i _02248_ _00551_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08593__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09051__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13035__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15639_ net1244 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XANTENNA__10197__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14892__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09160_ net979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[16\] net948 vssd1
+ vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09986__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08111_ _04519_ _04520_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17309_ clknet_leaf_127_wb_clk_i _02869_ _01172_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09091_ net992 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\] net945 vssd1
+ vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12616__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08042_ team_01_WB.instance_to_wrap.cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 _04473_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09006__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11349__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold901 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[6\] vssd1 vssd1 vccd1 vccd1
+ net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\] vssd1 vssd1 vccd1 vccd1
+ net2528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold934 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net2550
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold956 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold967 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[4\] net942 vssd1
+ vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12351__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1601 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net3217 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09226__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net3228 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11475__B _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[21\] net717 net683 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _08010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1634 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1 vccd1
+ net3250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13971__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1645 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net3261
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17616__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout640_A _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16059__A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1382_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08276__S net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09599__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\] net924 vssd1
+ vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__and3_1
XANTENNA__13026__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16640__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17766__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09896__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09358_ _05583_ _05620_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09245__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18193__1567 vssd1 vssd1 vccd1 vccd1 _18193__1567/HI net1567 sky130_fd_sc_hd__conb_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08309_ net1765 net2618 net1044 vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09289_ _05515_ _05551_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _06668_ _07582_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11251_ _05482_ _06982_ _07105_ _07185_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__a22o_1
XANTENNA__10273__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10202_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[1\] net957 vssd1
+ vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__A3 _07185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11182_ _06453_ net341 _07445_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10563__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[2\] net737 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__a22o_1
XANTENNA__12261__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15990_ net1327 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__inv_2
XANTENNA_input34_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ net1282 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
X_10064_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[3\] net927 vssd1
+ vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__and3_1
XANTENNA__08040__A team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17660_ clknet_leaf_15_wb_clk_i _03220_ _01523_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ net1340 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XANTENNA__08975__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17296__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ clknet_leaf_113_wb_clk_i _02239_ _00474_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13823_ team_01_WB.instance_to_wrap.cpu.c0.count\[9\] _04115_ vssd1 vssd1 vccd1 vccd1
+ _04116_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17591_ clknet_leaf_12_wb_clk_i _03151_ _01454_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13265__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10079__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16542_ clknet_leaf_64_wb_clk_i _02170_ _00405_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11276__C1 _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ _07718_ _04065_ net484 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__or3b_1
XFILLER_0_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ _05348_ _06922_ _06927_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__o31a_1
XANTENNA__09484__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ net2024 net199 net383 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08692__A0 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16473_ clknet_leaf_99_wb_clk_i _02101_ _00336_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09302__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ net772 _07456_ net968 vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a21oi_1
X_10897_ _05043_ _06807_ _05166_ _04988_ net509 net498 vssd1 vssd1 vccd1 vccd1 _07161_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18212_ net601 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15424_ net1275 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ net2499 net237 net391 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09236__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18143_ net1517 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15355_ net1317 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12567_ net2689 net209 net401 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__mux2_1
XANTENNA__12436__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14306_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\]
+ _04445_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ team_01_WB.instance_to_wrap.cpu.f0.i\[19\] _07758_ vssd1 vssd1 vccd1 vccd1
+ _07759_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18074_ net1448 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
X_15286_ net1303 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12498_ _08011_ _08012_ net488 vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__and3_2
Xhold208 _03316_ vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[6\] vssd1 vssd1 vccd1 vccd1
+ net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ clknet_leaf_135_wb_clk_i _02585_ _00888_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14237_ net793 _04232_ _04241_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__and3_1
X_11449_ _04618_ _07682_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10003__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ net1710 net585 _04327_ net1171 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[115\] net1727 net830 vssd1 vssd1
+ vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12171__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ net791 net790 _04236_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ clknet_leaf_108_wb_clk_i net2601 _01747_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1270 net1272 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__buf_4
Xfanout1281 net1284 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_4
X_08660_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[28\] net719 net713 vssd1
+ vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__a21o_1
X_17858_ clknet_leaf_78_wb_clk_i _03408_ _01678_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1292 net1301 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11046__A_N net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16809_ clknet_leaf_42_wb_clk_i _02369_ _00672_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13256__A0 team_01_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08591_ net1125 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\] net921
+ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and3_1
X_17789_ clknet_leaf_115_wb_clk_i _03347_ _01610_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16663__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11806__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09475__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _05472_ _05473_ _05474_ _05475_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__or4_1
XANTENNA__10358__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10490__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17019__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14220__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11034__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09143_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] net652 _05383_
+ _05392_ _05401_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12346__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08435__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A _07925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09074_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[18\] net626 _05322_ _05329_
+ _05333_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a2111o_1
X_18068__1442 vssd1 vssd1 vccd1 vccd1 _18068__1442/HI net1442 sky130_fd_sc_hd__conb_1
XFILLER_0_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17169__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1130_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold720 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[89\] vssd1 vssd1 vccd1 vccd1
+ net2347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10093__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1228_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold742 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\] vssd1 vssd1 vccd1 vccd1
+ net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 team_01_WB.instance_to_wrap.cpu.K0.enable vssd1 vssd1 vccd1 vccd1 net2369
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold775 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11742__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_A _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 _03463_ vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__A team_01_WB.instance_to_wrap.cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_1682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold797 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12081__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _06236_ _06237_ _06238_ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12298__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[21\] net646 _05171_
+ _05182_ _05183_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1420 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[20\] net847
+ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and3_1
Xhold1453 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net3080
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1475 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 net3091
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net3102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[27\] vssd1 vssd1 vccd1 vccd1
+ net3113 sky130_fd_sc_hd__dlygate4sd3_1
X_08789_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\] net656 net631 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a22o_1
X_10820_ net330 _06995_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10751_ _06414_ net505 vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__nor2_1
XANTENNA__08674__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09122__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10268__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13640__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13470_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _05550_ _05584_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__o211a_1
X_10682_ _04883_ _04905_ _06945_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14211__A2 _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net2331 net263 net420 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__mux2_1
XANTENNA__12256__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10565__A _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08977__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ net1269 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12352_ net2772 net271 net490 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
XANTENNA__08035__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10784__A1 _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11303_ net325 _07565_ _07566_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__or3b_1
X_15071_ net1293 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net2486 net216 net431 vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__mux2_1
XANTENNA__09926__B1 _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14022_ _04196_ _04197_ _04198_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__or3_2
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11234_ _05892_ _07496_ _06030_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11396__A _07121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11165_ _06524_ net339 net336 net511 _07428_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14278__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _06365_ _06370_ _06371_ _06372_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__nor4_1
X_15973_ net1334 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__inv_2
X_11096_ _05583_ net548 _05718_ _05923_ net503 net518 vssd1 vssd1 vccd1 vccd1 _07360_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[4\] net610 _06290_ _06295_
+ net673 vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__a2111o_1
X_17712_ clknet_leaf_110_wb_clk_i _03272_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14924_ net1251 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 team_01_WB.instance_to_wrap.cpu.f0.write_data\[2\] vssd1 vssd1 vccd1 vccd1
+ net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1
+ net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17643_ clknet_leaf_60_wb_clk_i _03203_ _01506_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14855_ net1354 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13806_ team_01_WB.instance_to_wrap.cpu.f0.i\[8\] team_01_WB.instance_to_wrap.cpu.f0.i\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17574_ clknet_leaf_141_wb_clk_i _03134_ _01437_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14786_ net1333 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11998_ net2916 net296 net468 vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16525_ clknet_leaf_61_wb_clk_i _02153_ _00388_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13737_ _04018_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08665__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ net534 _07208_ net546 vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ clknet_leaf_106_wb_clk_i _02084_ _00319_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_128_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09209__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13668_ _07986_ _03994_ net188 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__mux2_1
XANTENNA__09967__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14202__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15407_ net1251 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12619_ net2738 net263 net397 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16387_ clknet_leaf_84_wb_clk_i _00004_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13599_ _07931_ _03937_ net186 vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__mux2_1
X_18126_ net1500 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15338_ net1196 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18057_ net1433 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15269_ net1229 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13713__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17008_ clknet_leaf_23_wb_clk_i _02568_ _00871_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09917__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08196__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09830_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[7\] net893 vssd1
+ vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_2
Xfanout518 net519 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14269__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ _06020_ _06022_ _06024_ _05994_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18192__1566 vssd1 vssd1 vccd1 vccd1 _18192__1566/HI net1566 sky130_fd_sc_hd__conb_1
X_08712_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[23\] net715 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a22o_1
X_09692_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] net633 _05936_
+ _05939_ _05945_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_83_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ net578 _04902_ _04904_ _04883_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__o211a_1
XANTENNA__13229__A0 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_A _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[30\] net653 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08656__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1080_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout436_A _08022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10088__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1178_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12076__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1345_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ net1013 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] net865
+ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16559__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10766__A1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17804__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13696__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ net1002 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[18\] net872 vssd1
+ vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12804__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09908__B1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold550 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout972_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold583 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold594 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17954__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[5\] net870 vssd1
+ vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and3_1
XANTENNA__09117__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12970_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[4\] _07426_ net1035 vssd1 vssd1
+ vccd1 vccd1 _03654_ sky130_fd_sc_hd__mux2_1
XANTENNA__09687__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08956__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ net2555 net266 net477 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__mux2_1
Xhold1272 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12691__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1283 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11155__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14640_ net1401 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
X_11852_ net2863 net304 net479 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ net531 _07001_ _07060_ _07066_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14571_ net1409 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[21\] net676 net775 vssd1 vssd1
+ vccd1 vccd1 _07914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10454__A0 _06716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16310_ clknet_leaf_111_wb_clk_i _01944_ _00178_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13522_ net186 _03872_ _03873_ net771 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a211o_1
X_17290_ clknet_leaf_43_wb_clk_i _02850_ _01153_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ net533 _06995_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16241_ clknet_leaf_79_wb_clk_i _00021_ _00109_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13453_ _03804_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10665_ _06872_ _06878_ _06921_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12404_ net2983 net205 net421 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
X_16172_ clknet_leaf_58_wb_clk_i _01840_ _00040_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13384_ net2266 net329 net353 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1
+ vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10757__A1 _07020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ team_01_WB.instance_to_wrap.cpu.CU0.opcode\[5\] net764 vssd1 vssd1 vccd1
+ vccd1 _06860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ net1188 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12335_ net2671 net209 net492 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
XANTENNA__12714__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15054_ net1231 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12266_ _07842_ net495 _07845_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__and3_4
XANTENNA__10509__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14214__B net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__inv_2
X_11217_ _05890_ _06043_ _07370_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__nand3_1
XFILLER_0_120_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12197_ net2356 net294 net446 vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
XANTENNA__11704__A_N team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
X_11148_ _06598_ _06600_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09027__C net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15956_ net1330 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__inv_2
X_11079_ _07328_ _07329_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__o21a_1
X_18067__1441 vssd1 vssd1 vccd1 vccd1 _18067__1441/HI net1441 sky130_fd_sc_hd__conb_1
X_14907_ net1297 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15887_ net1353 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17626_ clknet_leaf_34_wb_clk_i _03186_ _01489_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14838_ net1343 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XANTENNA__10189__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14769_ net1177 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17557_ clknet_leaf_25_wb_clk_i _03117_ _01420_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10445__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ clknet_leaf_102_wb_clk_i net1890 _00371_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08290_ net3015 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[58\] net1050 vssd1 vssd1
+ vccd1 vccd1 _03457_ sky130_fd_sc_hd__mux2_1
X_17488_ clknet_leaf_24_wb_clk_i _03048_ _01351_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ clknet_leaf_77_wb_clk_i net2129 _00302_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09994__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11096__S1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ net1483 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12624__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17977__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14405__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08403__A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10652__B _05993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 _07970_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_2
Xfanout315 net317 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11173__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 _03750_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17207__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[7\] net905 vssd1
+ vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__and3_1
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout359 _03666_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_1
XANTENNA_fanout386_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] net846
+ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__and3_1
XANTENNA__09234__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] net879
+ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16231__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1295_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17357__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[29\] net625 net608 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[29\]
+ _04888_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08557_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\] net705 _04803_
+ _04808_ _04811_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout720_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__A0 _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout818_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12976__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10436__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08488_ net1108 net1111 net1114 net1106 vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and4b_1
XFILLER_0_33_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09841__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09400__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[26\] net658 net622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\]
+ _06713_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__a221o_1
XANTENNA__10739__A1 _06955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09109_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[17\] net739 net690 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a22o_1
XANTENNA__08801__A0 _05063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\] net649 net613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__a22o_1
XANTENNA__12534__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10843__A _06314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ net2314 net249 net453 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ net2412 net215 net459 vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold380 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[18\] vssd1 vssd1 vccd1 vccd1
+ net1996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10281__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _05138_ _06607_ _06610_ net344 vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12900__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10989__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 _04754_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08580__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout871 net874 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
X_15810_ net1307 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__inv_2
X_16790_ clknet_leaf_29_wb_clk_i _02350_ _00653_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout882 _04744_ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_4
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ net1283 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11393__B _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] net1055 net365 _03641_
+ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__a22o_1
XANTENNA__12664__A1 _07869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1080 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net3136 net238 net475 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15672_ net1242 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12884_ net1032 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1
+ vccd1 _03592_ sky130_fd_sc_hd__or2_2
XFILLER_0_34_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16724__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17411_ clknet_leaf_119_wb_clk_i _02971_ _01274_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14623_ net1372 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11835_ net780 _07954_ _07955_ _07956_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12709__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17342_ clknet_leaf_4_wb_clk_i _02902_ _01205_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08096__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ net1399 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XANTENNA__08096__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11766_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[24\] _07324_ net674 vssd1 vssd1
+ vccd1 vccd1 _07900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09832__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10737__B _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13505_ _03764_ _03766_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10717_ _06864_ _06865_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__nand2_1
X_17273_ clknet_leaf_125_wb_clk_i _02833_ _01136_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14485_ net1358 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11697_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__or2_1
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16224_ clknet_leaf_42_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[5\]
+ _00092_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ _03779_ _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09045__B1 _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18191__1565 vssd1 vssd1 vccd1 vccd1 _18191__1565/HI net1565 sky130_fd_sc_hd__conb_1
X_10648_ _05889_ _05852_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ net1331 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__inv_2
XANTENNA__11849__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ net2355 net329 net353 team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1
+ vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12444__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ _04799_ _06842_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__nand2_1
X_15106_ net1311 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
X_12318_ net2644 net248 net427 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
X_16086_ net1371 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__inv_2
X_13298_ net126 net808 net803 net1847 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ net1283 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12249_ net1783 net281 net437 vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09899__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16254__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08571__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16988_ clknet_leaf_14_wb_clk_i _02548_ _00851_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09054__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10115__C1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15939_ net1340 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09989__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ net996 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[12\] net856 vssd1
+ vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08411_ net1147 net1150 net1152 net1154 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__and4b_1
XFILLER_0_133_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17609_ clknet_leaf_38_wb_clk_i _03169_ _01472_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_09391_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[13\] net868
+ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__and3_1
XANTENNA__12619__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10418__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08342_ net2634 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[6\] net1041 vssd1 vssd1
+ vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
XANTENNA__13080__A1 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11091__B1 _07020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ net1791 net2138 net1050 vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09036__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12354__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_A _07984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1043_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11478__B _07701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09229__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08133__A _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1210_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1308_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13693__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout189 _07670_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08279__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _05985_ _05988_ _05989_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__or4_4
XANTENNA__12646__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09658_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] net708 net756 vssd1
+ vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08609_ _04869_ _04870_ _04871_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__or4_1
XANTENNA__12529__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[28\] net591 vssd1 vssd1 vccd1
+ vccd1 _05853_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11620_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[16\] net573 vssd1 vssd1 vccd1
+ vccd1 _07825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_132_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11551_ net1064 _07782_ _07783_ _07731_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09130__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10276__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\] net662 net623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14270_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[127\] _04233_ _04264_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[95\]
+ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__a221o_1
X_11482_ _04505_ _07699_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__nor2_2
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire557 _06025_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
XFILLER_0_80_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13221_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[21\]
+ net826 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
X_10433_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] net759 _06695_ _06696_
+ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__a22o_2
XANTENNA__12264__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18066__1440 vssd1 vssd1 vccd1 vccd1 _18066__1440/HI net1440 sky130_fd_sc_hd__conb_1
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10188__A2 _06450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input64_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ net2441 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[90\] net826 vssd1 vssd1
+ vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XANTENNA__09139__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[27\] net732 _04676_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[27\] _06616_ vssd1 vssd1 vccd1
+ vccd1 _06628_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ net3140 net191 net451 vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13083_ net558 _07807_ _03704_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__o21ai_1
X_17960_ clknet_leaf_100_wb_clk_i _03510_ _01780_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[0\] net667 _06543_ _06558_
+ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__o22a_4
XANTENNA__17522__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__A1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16911_ clknet_leaf_54_wb_clk_i _02471_ _00774_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12034_ net494 _08008_ _08012_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__and3_4
X_17891_ clknet_leaf_80_wb_clk_i _03441_ _01711_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12885__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12885__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16842_ clknet_leaf_43_wb_clk_i _02402_ _00705_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10896__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 _04691_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_8
XANTENNA__17672__CLK clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13985_ _03554_ _04163_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nand2_1
X_16773_ clknet_leaf_134_wb_clk_i _02333_ _00636_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12936_ net364 _03628_ _03629_ net1053 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__a32o_1
X_15724_ net1264 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XANTENNA__10112__A2 _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09602__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12867_ net1032 team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1
+ _03579_ sky130_fd_sc_hd__nor2_1
XANTENNA__12439__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15655_ net1184 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ net780 _07940_ _07941_ _07942_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__a2bb2o_4
X_14606_ net1378 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
X_15586_ net1290 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
X_12798_ net2254 net206 net373 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14537_ net1317 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
X_17325_ clknet_leaf_19_wb_clk_i _02885_ _01188_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11749_ net675 _07585_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ net1335 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
X_17256_ clknet_leaf_62_wb_clk_i _02816_ _01119_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ _03770_ _03771_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16207_ clknet_leaf_116_wb_clk_i _01874_ _00075_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_17187_ clknet_leaf_120_wb_clk_i _02747_ _01050_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12174__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14399_ net1310 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XANTENNA__10179__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11376__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16138_ net1322 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
XANTENNA__09049__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ net1133 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[19\] net962
+ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16069_ net1354 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13522__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08891_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[21\] net744 _05144_ _05145_
+ _05147_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14078__B1 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[9\] _04645_ net705 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09443_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[12\] net691 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10658__A _06919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12349__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_A _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ _05635_ _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13943__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14250__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08325_ net2358 net2626 net1046 vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout516_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10096__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1258_A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09009__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[92\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09885__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12084__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13356__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _04572_ _04581_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11367__A1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18021__1598 vssd1 vssd1 vccd1 vccd1 net1598 _18021__1598/LO sky130_fd_sc_hd__conb_1
XFILLER_0_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout885_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12812__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10080_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[3\] net703 _06331_ _06343_
+ net714 vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18190__1564 vssd1 vssd1 vccd1 vccd1 _18190__1564/HI net1564 sky130_fd_sc_hd__conb_1
XFILLER_0_96_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13770_ net1662 net782 _04078_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10982_ _05482_ _07244_ _05419_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ net2080 net244 net385 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15440_ net1256 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net2830 net262 net392 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17075__CLK clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09248__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A team_01_WB.instance_to_wrap.cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14241__B1 _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ net496 _07816_ net3213 net838 vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o2bb2a_1
X_15371_ net1210 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XANTENNA__13595__A2 _07243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ net2860 net247 net399 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17110_ clknet_leaf_29_wb_clk_i _02670_ _00973_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14322_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\]
+ _04455_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__and3_1
X_18090_ net1464 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
X_11534_ team_01_WB.instance_to_wrap.cpu.f0.i\[4\] net1161 _07722_ vssd1 vssd1 vccd1
+ vccd1 _07769_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17041_ clknet_leaf_20_wb_clk_i _02601_ _00904_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14253_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[78\] _04246_ _04263_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[70\]
+ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a22o_1
X_11465_ _04468_ _07717_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13204_ net3061 net2820 net819 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XANTENNA__13752__C1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ net970 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[26\] net935 vssd1
+ vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__and3_1
X_14184_ _04244_ _04276_ _04340_ _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11396_ _07121_ _07152_ _07653_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__and3_1
XANTENNA__16912__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13135_ net1767 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\] net831 vssd1 vssd1
+ vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XANTENNA__12722__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10347_ _05211_ _06610_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13066_ _05414_ _07803_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__nand2_1
X_17943_ clknet_leaf_109_wb_clk_i net3003 _01763_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[0\] net636 _06539_ _06540_
+ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__a2111o_1
X_12017_ net2165 net280 net464 vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XANTENNA__08526__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17874_ clknet_leaf_78_wb_clk_i _03424_ _01694_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16825_ clknet_leaf_125_wb_clk_i _02385_ _00688_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13553__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13283__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16756_ clknet_leaf_7_wb_clk_i _02316_ _00619_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13968_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[1\] net584 vssd1 vssd1
+ vccd1 vccd1 _04161_ sky130_fd_sc_hd__or2_1
XANTENNA__09332__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15707_ net1317 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
X_12919_ net3258 net604 net586 _03617_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12169__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16687_ clknet_leaf_93_wb_clk_i _02247_ _00550_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13899_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[12\] net795 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[12\] sky130_fd_sc_hd__and2_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15638_ net1304 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09239__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14232__B1 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16442__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15569_ net1200 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17568__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ _04515_ _04516_ _04521_ _04522_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17308_ clknet_leaf_10_wb_clk_i _02868_ _01171_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09090_ net983 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\] _04657_
+ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08041_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1 _04472_
+ sky130_fd_sc_hd__inv_2
X_17239_ clknet_leaf_9_wb_clk_i _02799_ _01102_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11102__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold902 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold913 _02128_ vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold935 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold946 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold957 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 team_01_WB.instance_to_wrap.cpu.f0.num\[11\] vssd1 vssd1 vccd1 vccd1 net2584
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15509__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ net989 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[4\] net942 vssd1
+ vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
XANTENNA__12632__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold979 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14413__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08943_ _05070_ _05138_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__nor3_1
XANTENNA__10660__B _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout299_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08517__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1602 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 net3218
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08874_ _05136_ _05137_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or2_2
Xhold1613 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net3229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1006_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1624 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1635 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3251 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1646 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net3262
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17098__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09478__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__B2 team_01_WB.instance_to_wrap.a1.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08784__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12079__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09426_ net972 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[12\] net950 vssd1
+ vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14223__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13699__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09357_ _05583_ _05620_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12807__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08308_ net2061 net3120 net1039 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ _05515_ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08239_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[117\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[109\]
+ net1042 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13734__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net331 _05484_ _05481_ net335 vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10201_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] net915 vssd1
+ vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08756__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ _06453_ net339 net336 net530 net333 vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__a221o_1
XANTENNA__12542__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08959__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[2\] net932 vssd1
+ vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14940_ net1234 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
X_10063_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[3\] net939 vssd1
+ vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10315__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ net1340 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16610_ clknet_leaf_112_wb_clk_i _02238_ _00473_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15154__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13822_ team_01_WB.instance_to_wrap.cpu.c0.count\[8\] team_01_WB.instance_to_wrap.cpu.c0.count\[7\]
+ _04113_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17590_ clknet_leaf_29_wb_clk_i _03150_ _01453_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16541_ clknet_leaf_64_wb_clk_i _02169_ _00404_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13753_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] _07716_ vssd1 vssd1 vccd1 vccd1
+ _04065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11276__B1 _06867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10965_ net323 _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12704_ net2390 net288 net383 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
XANTENNA__17710__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13684_ net770 _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nand2_1
X_16472_ clknet_leaf_106_wb_clk_i _02100_ _00335_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10896_ _05205_ _06873_ _07158_ net322 vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18211_ net1585 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
X_15423_ net1295 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
X_12635_ net2987 net205 net393 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12717__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11579__A1 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13402__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18142_ net1516 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
XFILLER_0_81_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15354_ net1305 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ net2462 net192 net399 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17860__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ _07701_ _07757_ net319 vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14305_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] _04445_ net1830 vssd1
+ vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18073_ net1447 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
X_15285_ net1173 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
X_12497_ net2234 net213 net414 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold209 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ _04345_ _04392_ _04373_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__a21oi_1
X_17024_ clknet_leaf_141_wb_clk_i _02584_ _00887_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11448_ _04618_ _07682_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__nor2_4
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14167_ _04319_ _04324_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or4_1
XANTENNA__12452__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _06937_ net322 _07127_ _07642_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13118_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[124\]
+ net818 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ net793 net790 net787 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[23\] _03685_ net1028 vssd1
+ vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ clknet_leaf_101_wb_clk_i _03476_ _01746_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_98_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__buf_4
XANTENNA__17240__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1271 net1272 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_2
Xfanout1282 net1284 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ clknet_leaf_106_wb_clk_i _03407_ _01677_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1293 net1296 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_4
XFILLER_0_117_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15064__A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16808_ clknet_leaf_45_wb_clk_i _02368_ _00671_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16808__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ _04852_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17788_ clknet_leaf_114_wb_clk_i _03346_ _01609_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15999__A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16739_ clknet_leaf_131_wb_clk_i _02299_ _00602_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11806__A2 _07265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18020__1597 vssd1 vssd1 vccd1 vccd1 net1597 _18020__1597/LO sky130_fd_sc_hd__conb_1
XFILLER_0_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09997__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14205__B1 _04244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[16\] net656 _05457_
+ _05460_ _05464_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16958__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12627__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09142_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[17\] net621 _05387_
+ _05388_ _05397_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] net624 _05321_ _05324_
+ _05326_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout214_A _08007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold710 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold721 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold743 _03430_ vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12362__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold754 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 net2370
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold765 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10545__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09975_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[5\] net649 _06215_ _06219_
+ _06220_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__a2111o_1
Xhold798 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08926_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[21\] net608 _05172_
+ _05176_ _05184_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__a2111o_1
Xhold1410 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net3026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net3037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[107\] vssd1 vssd1 vccd1 vccd1
+ net3048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[20\] net849
+ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__and3_1
Xhold1443 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net3059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout750_A _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1454 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3070 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16488__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1465 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[8\] vssd1 vssd1 vccd1 vccd1
+ net3081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1476 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1487 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3103 sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ _05045_ _05047_ _05049_ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nor4_1
Xhold1498 _03426_ vssd1 vssd1 vccd1 vccd1 net3114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09403__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _07012_ _07013_ net517 vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09700__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\] net638 net626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17883__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ _06840_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__nor2_1
XANTENNA__12537__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10218__D1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ net2595 net266 net421 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12351_ net2567 net247 net491 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11302_ _05962_ _07552_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__nand2_1
X_15070_ net1297 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ net2018 net279 net432 vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[14\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[17\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__or4bb_1
X_11233_ _05892_ _06030_ _07496_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__and3_1
XANTENNA__12272__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__A team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11733__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11164_ _06485_ net511 net333 vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o21a_1
XANTENNA__17263__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\] net641 _06378_ net673
+ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_78_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15972_ net1334 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__inv_2
X_11095_ _05718_ _05923_ net503 vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__mux2_1
XANTENNA__08986__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ clknet_leaf_110_wb_clk_i _03271_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ _06306_ _06307_ _06308_ _06309_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__or4_2
X_14923_ net1208 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold70 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1 vccd1
+ net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_01_WB.instance_to_wrap.cpu.f0.write_data\[27\] vssd1 vssd1 vccd1 vccd1
+ net1697 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ clknet_leaf_41_wb_clk_i _03202_ _01505_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold92 team_01_WB.instance_to_wrap.cpu.f0.read_i vssd1 vssd1 vccd1 vccd1 net1708
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08901__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__A1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14854_ net1354 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13805_ net1673 net784 _04105_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__o21a_1
XANTENNA__13789__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17573_ clknet_leaf_135_wb_clk_i _03133_ _01436_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11997_ net2723 net307 net468 vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
X_14785_ net1387 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16524_ clknet_leaf_59_wb_clk_i _02152_ _00387_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13736_ net1062 _04017_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__nand2_1
X_10948_ net540 _07211_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__nand2_1
XANTENNA__09862__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09610__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16455_ clknet_leaf_81_wb_clk_i _02083_ _00318_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13667_ _03778_ _03790_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879_ _07029_ _07049_ net522 vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__mux2_1
XANTENNA__12447__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15406_ net1229 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12618_ net3223 net268 net397 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
X_16386_ clknet_leaf_84_wb_clk_i _00003_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13598_ _03832_ _03936_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08968__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18125_ net1499 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
X_15337_ net1214 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
X_12549_ net2192 net274 net404 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__mux2_1
XANTENNA__10194__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_1 _07962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18056_ net1432 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_124_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15268_ net1270 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
XANTENNA__17606__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17007_ clknet_leaf_18_wb_clk_i _02567_ _00870_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14219_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\] _04229_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\]
+ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__a22o_1
XANTENNA__12182__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15199_ net1293 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10527__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout508 _06560_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_2
Xfanout519 _06522_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09760_ _06013_ _06014_ _06015_ _06023_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__or4_1
XANTENNA__16630__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] net721 _04961_
+ _04962_ _04973_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11488__B1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17909_ clknet_leaf_104_wb_clk_i _03459_ _01729_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[68\]
+ sky130_fd_sc_hd__dfstp_1
X_09691_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[11\] net612 _05937_ _05943_
+ _05944_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
X_08642_ _04883_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08573_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\] net628 _04836_
+ net670 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11660__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout331_A _06989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12357__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout429_A _08024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09125_ net1075 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[17\] net865
+ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__and3_1
XANTENNA__13977__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09081__A1 _05344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1240_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1338_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[18\] net872
+ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16160__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17286__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09893__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13188__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 net2156
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12092__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold551 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold562 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[26\] vssd1 vssd1 vccd1 vccd1
+ net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold573 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09384__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold584 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold595 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12820__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14601__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ net1089 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] net908 vssd1
+ vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08909_ net1012 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[21\] net879
+ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09889_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[6\] net883 vssd1
+ vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 _03509_ vssd1 vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[50\] vssd1 vssd1 vccd1 vccd1
+ net2867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1262 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ net2520 net270 net475 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__mux2_1
Xhold1273 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ net2889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1284 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11851_ _07968_ _07969_ net780 vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__mux2_4
XANTENNA__09133__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13651__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ net531 _07050_ _07065_ net321 vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__o211a_1
XANTENNA__15432__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14570_ net1355 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ net676 _07196_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09430__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13521_ net185 _07871_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__nor2_1
X_10733_ net538 _06996_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11651__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ clknet_leaf_90_wb_clk_i _00020_ _00108_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13452_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] net592 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a21oi_1
X_10664_ _05281_ _06924_ _06927_ _06878_ _06923_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__a221o_1
XANTENNA__14196__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16503__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08046__A team_01_WB.instance_to_wrap.cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12403_ net2857 net238 net419 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13383_ net3101 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[15\] vssd1 vssd1
+ vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
X_16171_ clknet_leaf_58_wb_clk_i _01839_ _00039_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10595_ team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] _06851_ vssd1 vssd1 vccd1
+ vccd1 _06859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ net2836 net192 net490 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
X_15122_ net1178 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13098__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15053_ net1216 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
X_12265_ net3235 net210 net438 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17779__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16653__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14004_ _03555_ _04181_ _03556_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12903__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11216_ _07379_ _07396_ _07414_ _07479_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__and4b_1
XANTENNA__09375__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net2620 net307 net446 vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
XANTENNA__11182__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11147_ _06972_ _07183_ _07399_ _07402_ _07410_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__o2111a_1
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__12730__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10390__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17009__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14120__A2 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15955_ net1330 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__inv_2
X_11078_ _07107_ _07340_ _07341_ _07332_ _07338_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__o311a_1
X_10029_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[4\] net852 vssd1
+ vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__and3_1
X_14906_ net1306 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
X_15886_ net1357 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17625_ clknet_leaf_16_wb_clk_i _03185_ _01488_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14837_ net1343 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11870__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08638__A1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[29\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17556_ clknet_leaf_4_wb_clk_i _03116_ _01419_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ net1237 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08882__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16507_ clknet_leaf_101_wb_clk_i net3130 _00370_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ _04028_ _04038_ net485 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12177__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17487_ clknet_leaf_124_wb_clk_i _03047_ _01350_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14699_ net1363 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14187__A2 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16438_ clknet_leaf_80_wb_clk_i _02066_ _00301_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16183__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16369_ clknet_leaf_66_wb_clk_i net1828 _00237_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11945__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18108_ net1482 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18039_ net1429 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_1_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08403__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _07970_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_2
XANTENNA__08574__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout327 _03750_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09812_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[7\] net887 vssd1
+ vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__and3_1
XANTENNA__12640__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout338 _06983_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_4
Xfanout349 _04569_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10381__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09743_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[10\] net861
+ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout281_A _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout379_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ net1024 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\] net883 vssd1
+ vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10133__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08625_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] net661 net649 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1190_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08556_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\] net691 _04804_
+ _04805_ _04809_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09888__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ net1001 net867 vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__and2_2
XANTENNA__12087__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout713_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14178__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12189__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12815__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[17\] net704 net696 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[17\]
+ _05350_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a221o_1
XANTENNA__17921__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10380_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[27\] net657 net615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09039_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[18\] net749 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[18\]
+ _05289_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12050_ net2169 net278 net461 vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
Xhold370 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold381 net106 vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09128__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11001_ net346 _07245_ _07246_ _07264_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__a31o_2
Xhold392 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12550__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10372__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net854 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 _04754_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_2
XANTENNA__09109__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout872 net874 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout883 net884 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_4
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_4
X_15740_ net1278 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
X_12952_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[9\] _07495_ net1034 vssd1 vssd1
+ vccd1 vccd1 _03641_ sky130_fd_sc_hd__mux2_1
Xhold1070 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\] vssd1 vssd1 vccd1 vccd1
+ net2686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1081 team_01_WB.instance_to_wrap.cpu.f0.num\[10\] vssd1 vssd1 vccd1 vccd1 net2697
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11903_ net2530 net206 net477 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__mux2_1
Xhold1092 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15671_ net1238 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
X_12883_ net1025 _07640_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17410_ clknet_leaf_143_wb_clk_i _02970_ _01273_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14622_ net1378 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11834_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[12\] net679 net776 vssd1 vssd1
+ vccd1 vccd1 _07956_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17341_ clknet_leaf_127_wb_clk_i _02901_ _01204_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14553_ net1407 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
X_11765_ net774 _07898_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_82_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13504_ _03767_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ _06866_ _06978_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14169__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17272_ clknet_leaf_28_wb_clk_i _02832_ _01135_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11696_ net2909 net153 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03257_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14484_ net1385 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16223_ clknet_leaf_42_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[4\]
+ _00091_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09045__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13435_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[4\] _06278_ vssd1 vssd1 vccd1
+ vccd1 _03788_ sky130_fd_sc_hd__or2_1
X_10647_ _06036_ _06910_ _06909_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__a21o_1
XANTENNA__12725__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ net1332 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__inv_2
X_13366_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _03749_ vssd1 vssd1 vccd1 vccd1
+ _03751_ sky130_fd_sc_hd__nor2_1
X_10578_ _04853_ _06841_ _04852_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__a21o_1
XANTENNA__08504__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ net1291 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12317_ net1825 net275 net428 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
X_13297_ net127 net810 net805 net1694 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
X_16085_ net1348 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__inv_2
XANTENNA__08223__B _04617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__C net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15036_ net1280 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
X_12248_ net3029 net252 net436 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11865__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15337__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ net1982 net282 net443 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__mux2_1
XANTENNA__10363__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08877__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ clknet_leaf_37_wb_clk_i _02547_ _00850_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_15938_ net1308 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16549__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15869_ net1393 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08410_ net974 net929 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__and2_2
X_17608_ clknet_leaf_46_wb_clk_i _03168_ _01471_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15072__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] net669 vssd1 vssd1
+ vccd1 vccd1 _05654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08341_ net2710 net2965 net1044 vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__mux2_1
X_17539_ clknet_leaf_120_wb_clk_i _03099_ _01402_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09501__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16699__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13080__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[76\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
XANTENNA__17944__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__B2 _06971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18159__1533 vssd1 vssd1 vccd1 vccd1 _18159__1533/HI net1533 sky130_fd_sc_hd__conb_1
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12635__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08414__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08795__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1036_A team_01_WB.instance_to_wrap.cpu.RU0.InstrRead vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13974__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13540__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12370__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13693__C team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18115__1489 vssd1 vssd1 vccd1 vccd1 _18115__1489/HI net1489 sky130_fd_sc_hd__conb_1
XFILLER_0_138_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout663_A _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[10\] net733 net724 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[10\]
+ _05979_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09511__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ net713 _05911_ _05916_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout928_A _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[29\] net747 _04861_
+ _04862_ _04866_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a2111o_1
X_09588_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[8\] net761 _05850_ _05851_
+ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a22o_2
XANTENNA__08295__S net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08539_ net1119 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\] net929
+ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11550_ net1064 _07781_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__nor2_1
XANTENNA__15710__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[25\] net647 _06762_
+ _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13359__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11481_ _07733_ _07730_ team_01_WB.instance_to_wrap.cpu.f0.i\[31\] vssd1 vssd1 vccd1
+ vccd1 _03379_ sky130_fd_sc_hd__mux2_1
XANTENNA__12545__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ net2568 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[22\] net820 vssd1 vssd1
+ vccd1 vccd1 _02038_ sky130_fd_sc_hd__mux2_1
Xwire558 _05751_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_4
XANTENNA__09578__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[26\] net707 net755 vssd1
+ vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08786__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\] net2455 net830 vssd1 vssd1
+ vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[27\] net752 net699 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10292__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ net2290 net196 net452 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
X_13082_ net356 _03707_ _03708_ net835 net3156 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a32o_1
X_10294_ _06547_ _06549_ _06553_ _06557_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__or4_1
XANTENNA_input57_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12033_ net3014 net214 net465 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
X_16910_ clknet_leaf_52_wb_clk_i _02470_ _00773_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12280__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17890_ clknet_leaf_75_wb_clk_i net3053 _01710_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08697__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09155__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16841_ clknet_leaf_41_wb_clk_i _02401_ _00704_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09750__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _04718_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout691 net694 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_16772_ clknet_leaf_128_wb_clk_i _02332_ _00635_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ _03558_ _04171_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__and2_1
X_15723_ net1208 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
X_12935_ net1030 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1
+ vccd1 _03629_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11845__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219__1587 vssd1 vssd1 vccd1 vccd1 _18219__1587/HI net1587 sky130_fd_sc_hd__conb_1
XANTENNA__08710__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16841__CLK clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13405__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15654_ net1275 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XANTENNA__17967__CLK clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12866_ team_01_WB.instance_to_wrap.cpu.DM0.state\[0\] _07834_ team_01_WB.instance_to_wrap.cpu.DM0.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14605_ net1375 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
X_11817_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[15\] net676 net776 vssd1 vssd1
+ vccd1 vccd1 _07942_ sky130_fd_sc_hd__o21a_1
XANTENNA__09321__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15585_ net1313 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12797_ net2418 net192 net371 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10467__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ clknet_leaf_44_wb_clk_i _02884_ _01187_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14536_ net1318 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[27\] _07863_ vssd1 vssd1
+ vccd1 vccd1 _07885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ clknet_leaf_131_wb_clk_i _02815_ _01118_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14467_ net1336 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
XANTENNA__12455__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ net1651 net1160 net568 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16206_ clknet_leaf_116_wb_clk_i _01873_ _00074_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13418_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] net591 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17186_ clknet_leaf_0_wb_clk_i _02746_ _01049_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14398_ net1310 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16137_ net1321 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ net7 net801 net596 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\] vssd1 vssd1
+ vccd1 vccd1 _01931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16068_ net1403 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09991__C net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08529__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15019_ net1205 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XANTENNA__12190__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08890_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[21\] net726 net713 _05140_
+ _05143_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09065__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__A_N net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09511_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[9\] net753 _04680_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08701__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ _05703_ _05704_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__or3_1
XANTENNA__08409__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13589__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[13\] net731 net715 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a22o_1
XANTENNA__09231__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13053__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08128__B _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08324_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\] net2504 net1039 vssd1 vssd1
+ vccd1 vccd1 _03423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08255_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[93\]
+ net1043 vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XANTENNA__14146__A _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout411_A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout509_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1153_A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08186_ _04571_ _04581_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08768__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1261_A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout878_A _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10327__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09406__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16864__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13816__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09703__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[10\] net937
+ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and3_1
X_10981_ _05419_ _05482_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ net2938 net315 net384 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ net2127 net267 net393 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10287__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[25\] net572 vssd1 vssd1 vccd1
+ vccd1 _07816_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ net2200 net274 net400 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__mux2_1
X_15370_ net1201 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14321_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[15\] _04455_ net1780 vssd1
+ vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a21oi_1
X_11533_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] _07745_ _07766_ _07768_ vssd1
+ vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o211a_1
XANTENNA__16244__CLK clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12275__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08471__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ clknet_leaf_23_wb_clk_i _02600_ _00903_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11464_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__inv_2
X_14252_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\] _04272_ _04276_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[46\]
+ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10415_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\] net920
+ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and3_1
X_13203_ net2617 net1732 net825 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
X_14183_ _04252_ _04253_ _04269_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__or4_1
X_11395_ _07223_ _07522_ _07656_ _07658_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16394__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13134_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[100\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[108\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
X_10346_ _05279_ _06609_ _06608_ _05349_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_123_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09971__A2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ net1712 net835 net356 _03696_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
X_17942_ clknet_leaf_103_wb_clk_i _03492_ _01762_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[101\]
+ sky130_fd_sc_hd__dfstp_1
X_10277_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\] net859 vssd1
+ vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08501__B net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09184__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ net2404 net253 net465 vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
XANTENNA__09723__A2 _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17873_ clknet_leaf_109_wb_clk_i net2505 _01693_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_18158__1532 vssd1 vssd1 vccd1 vccd1 _18158__1532/HI net1532 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16824_ clknet_leaf_28_wb_clk_i _02384_ _00687_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12958__B _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16755_ clknet_leaf_48_wb_clk_i _02315_ _00618_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__inv_2
XANTENNA__13283__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ net1259 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
X_12918_ net364 _03615_ _03616_ net1054 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__a32o_1
X_16686_ clknet_leaf_55_wb_clk_i _02246_ _00549_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] net797 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[11\] sky130_fd_sc_hd__and2_1
X_15637_ net1179 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09051__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ net2186 net266 net369 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10197__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ net1250 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XANTENNA__09986__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17307_ clknet_leaf_36_wb_clk_i _02867_ _01170_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10254__C1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14519_ net1411 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12185__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18114__1488 vssd1 vssd1 vccd1 vccd1 _18114__1488/HI net1488 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ net1211 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08040_ team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _04471_
+ sky130_fd_sc_hd__inv_2
X_17238_ clknet_leaf_33_wb_clk_i _02798_ _01101_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16737__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12546__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold903 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11102__B _07365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17169_ clknet_leaf_22_wb_clk_i _02729_ _01032_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold914 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10557__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[22\] vssd1 vssd1 vccd1 vccd1
+ net2552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold947 team_01_WB.instance_to_wrap.cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1 net2563
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold958 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net1144 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] net959 vssd1
+ vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__and3_1
Xhold969 _01896_ vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08942_ _05203_ _05204_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__or2_2
XANTENNA__16887__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _05099_ _05135_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nor2_1
Xhold1603 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09226__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1614 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3230 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1625 team_01_WB.instance_to_wrap.cpu.SR1.char_in\[4\] vssd1 vssd1 vccd1 vccd1
+ net3241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1636 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1647 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 net3263
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11809__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout361_A _03665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout459_A _08015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11285__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08150__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09425_ net548 _05687_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16267__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1270_A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout626_A _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1368_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ net582 net559 _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09896__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_139_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11588__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[49\] net3052 net1048 vssd1 vssd1
+ vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XANTENNA__12095__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ _05549_ _05550_ net580 vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08238_ net2855 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[110\] net1039 vssd1 vssd1
+ vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17662__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout995_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08169_ team_01_WB.instance_to_wrap.cpu.K0.code\[7\] team_01_WB.instance_to_wrap.cpu.K0.code\[5\]
+ team_01_WB.instance_to_wrap.cpu.K0.code\[4\] team_01_WB.instance_to_wrap.cpu.K0.code\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or4b_2
XANTENNA__12823__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10548__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[1\] net928 vssd1
+ vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11180_ _06456_ _06883_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08602__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10131_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[2\] _04655_ vssd1
+ vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10062_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] net959 vssd1
+ vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__and3_1
XANTENNA__09136__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14870_ net1345 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17042__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ team_01_WB.instance_to_wrap.cpu.c0.count\[7\] _04113_ vssd1 vssd1 vccd1 vccd1
+ _04114_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09433__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13265__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10079__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16540_ clknet_leaf_56_wb_clk_i _02168_ _00403_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13752_ _07718_ _07773_ _04016_ _04468_ _04558_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a221o_1
X_10964_ _06922_ _06927_ _05348_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__o21a_1
XANTENNA__08049__A team_01_WB.instance_to_wrap.cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12703_ net2468 net231 net385 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
X_16471_ clknet_leaf_76_wb_clk_i net2749 _00334_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_13683_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] _04006_ net187 vssd1
+ vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__mux2_1
X_10895_ _05138_ _05206_ _07157_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11902__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18210_ net1584 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
X_15422_ net1291 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ net2708 net240 net393 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18141_ net1515 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
XFILLER_0_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11123__S1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15353_ net1192 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10787__A0 _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08444__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ net2224 net195 net401 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304_ net3025 _04445_ _04447_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__o21a_1
XANTENNA__10251__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ _07714_ _07739_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__and2_1
X_18072_ net1446 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15284_ net1240 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12496_ net1943 net290 net412 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ clknet_leaf_3_wb_clk_i _02583_ _00886_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14235_ _04382_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nor2_1
X_11447_ _04560_ _07699_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__or2_1
XANTENNA__12733__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09947__A1_N _06209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14166_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[10\] _04267_ _04288_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ _04158_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a221o_1
X_11378_ _06778_ _06936_ _07126_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output88_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08512__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ net505 _06591_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13117_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\]
+ net823 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ net791 net788 _04237_ _04258_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[88\]
+ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14150__B1 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13933__A_N net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ _05009_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ clknet_leaf_105_wb_clk_i _03475_ _01745_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[84\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1250 net1253 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_4
Xfanout1261 net1268 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17856_ clknet_leaf_99_wb_clk_i _03406_ _01676_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1272 net1301 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__clkbuf_4
Xfanout1283 net1284 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_2
Xfanout1294 net1296 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__buf_4
XANTENNA__09343__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ clknet_leaf_130_wb_clk_i _02367_ _00670_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08885__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17787_ clknet_leaf_113_wb_clk_i _03345_ _01608_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10489__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14999_ net1244 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17535__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16738_ clknet_leaf_142_wb_clk_i _02298_ _00601_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16669_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[23\]
+ _00532_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08683__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[16\] net626 _05453_ _05459_
+ _05466_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09489__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10490__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12767__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[17\] net619 _05395_
+ _05398_ _05400_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08435__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09072_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[18\] net631 _05323_
+ _05327_ _05332_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12643__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold700 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold711 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A _07879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold722 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[17\] vssd1 vssd1 vccd1 vccd1
+ net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 team_01_WB.instance_to_wrap.cpu.f0.write_data\[26\] vssd1 vssd1 vccd1 vccd1
+ net2349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold744 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08422__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold766 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 net2382
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold777 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[5\] net643 _06214_ _06227_
+ _06231_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a2111o_1
Xhold799 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\] vssd1 vssd1 vccd1 vccd1
+ net2415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08141__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17065__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14141__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[21\] net635 net620 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1400 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1411 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _02131_ vssd1 vssd1 vccd1 vccd1 net3049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08856_ net999 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[20\] net877 vssd1
+ vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__and3_1
Xhold1444 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net3060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net3071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net3082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1477 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 net3093
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout743_A _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[22\] net646 net612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[22\]
+ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a221o_1
Xhold1488 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net3104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1499 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout910_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08674__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[13\] net860
+ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10481__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ _04956_ _04935_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_113_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ net1001 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[14\] net909 vssd1
+ vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18157__1531 vssd1 vssd1 vccd1 vccd1 _18157__1531/HI net1531 sky130_fd_sc_hd__conb_1
X_12350_ net2969 net276 net491 vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11301_ _05962_ _07552_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12281_ net1950 net252 net433 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__mux2_1
XANTENNA__12553__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14334__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14020_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[13\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[12\]
+ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[11\] team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09387__B1 _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ _06602_ _06603_ _06041_ _06043_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__a211o_1
XANTENNA__09926__A2 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11163_ _06996_ _07252_ _07261_ net330 vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11396__C _07653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14132__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] net665 net623 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ net1332 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__inv_2
X_11094_ _07356_ _07357_ net517 vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__mux2_1
X_17710_ clknet_leaf_109_wb_clk_i _03270_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16432__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[4\] net654 _06284_ _06287_
+ _06291_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17558__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14922_ net1197 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18113__1487 vssd1 vssd1 vccd1 vccd1 _18113__1487/HI net1487 sky130_fd_sc_hd__conb_1
Xhold60 net151 vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_01_WB.instance_to_wrap.cpu.f0.write_data\[12\] vssd1 vssd1 vccd1 vccd1
+ net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 net138 vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ clknet_leaf_22_wb_clk_i _03201_ _01504_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09163__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14853_ net1350 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
Xhold93 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[5\] vssd1 vssd1 vccd1 vccd1
+ net1709 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ _04556_ _07704_ _04102_ _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__a31o_1
X_17572_ clknet_leaf_138_wb_clk_i _03132_ _01435_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14784_ net1399 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
X_11996_ net2783 net312 net468 vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08114__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16523_ clknet_leaf_75_wb_clk_i _02151_ _00386_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13735_ team_01_WB.instance_to_wrap.cpu.f0.data_adr\[26\] net782 _04051_ vssd1 vssd1
+ vccd1 vccd1 _01848_ sky130_fd_sc_hd__o21a_1
XANTENNA__12728__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10947_ _07209_ _07210_ net525 vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08665__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13413__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14199__B1 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16454_ clknet_leaf_80_wb_clk_i _02082_ _00317_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13666_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[6\] _03993_ net1067 vssd1
+ vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XANTENNA__08507__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ _06998_ _07133_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15405_ net1215 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12617_ net2912 net272 net395 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
X_16385_ clknet_leaf_83_wb_clk_i _00002_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13597_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] _05449_ _03829_ vssd1
+ vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18124_ net1498 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
XFILLER_0_14_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15336_ net1204 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
X_12548_ net1989 net217 net403 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18055_ net1431 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__12463__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15267_ net1225 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
X_12479_ net2111 net254 net412 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17006_ clknet_leaf_52_wb_clk_i _02566_ _00869_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09378__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17088__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\] _04227_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[85\]
+ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09917__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15198_ net1315 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12921__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[66\] _04272_ _04273_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__a22o_1
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08710_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\] net725 net701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a22o_1
X_17908_ clknet_leaf_76_wb_clk_i _03458_ _01728_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_09690_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\] net663 _05927_
+ _05929_ _05932_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_83_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1080 net1096 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_2
X_08641_ net578 _04902_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o21ai_1
XANTENNA__16925__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1091 net1096 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_2
X_17839_ clknet_leaf_84_wb_clk_i _03390_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08572_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[30\] net644 net616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09838__D1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12638__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08656__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11660__B2 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08417__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\] net893 vssd1
+ vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__and3_1
XANTENNA__16305__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09055_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[18\] net863
+ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12373__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11497__B _07734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1 vccd1
+ net2146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09908__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold541 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold552 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[19\] vssd1 vssd1 vccd1 vccd1
+ net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1400_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold596 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[5\] net879 vssd1
+ vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout860_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout958_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08908_ net1014 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] net893 vssd1
+ vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__and3_1
X_09888_ net1099 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[6\] net858 vssd1
+ vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__and3_1
Xhold1230 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1241 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ net1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[20\] net908
+ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__and3_1
XANTENNA__17850__CLK clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1263 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__A1 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1274 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\] vssd1 vssd1 vccd1 vccd1
+ net2890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__B2 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1285 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15713__A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1296 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11850_ team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\] _07495_ net679 vssd1 vssd1
+ vccd1 vccd1 _07969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12979__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ net527 _07053_ _07062_ _07064_ net537 vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12979__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11781_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[21\] _07859_ vssd1 vssd1
+ vccd1 vccd1 _07912_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12548__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _03754_ _03866_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10732_ _06952_ _06978_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11651__B2 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[29\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\]
+ net592 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10663_ _05378_ _05415_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12402_ net1994 net208 net421 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__mux2_1
XANTENNA__10206__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16170_ clknet_leaf_57_wb_clk_i _01838_ _00038_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13382_ net2410 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[16\] vssd1 vssd1
+ vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10594_ _04632_ _06846_ _06847_ _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09072__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15121_ net1199 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12333_ net2759 net195 net492 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12283__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15052_ net1263 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
X_12264_ net2777 net291 net437 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11167__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14003_ _04164_ _03553_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__or2_1
XANTENNA__12903__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11215_ _07426_ _07441_ _07456_ _07478_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__and4b_1
XANTENNA__12903__B2 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12195_ net3149 net312 net446 vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17380__CLK clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08583__B2 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16948__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11146_ _07106_ _07409_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13408__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15954_ net1330 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__inv_2
X_11077_ net536 _07272_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10028_ net1094 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[4\] net869 vssd1
+ vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__and3_1
X_14905_ net1244 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09324__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15885_ net1359 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17624_ clknet_leaf_27_wb_clk_i _03184_ _01487_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14836_ net1343 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XANTENNA__12966__B _07414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17555_ clknet_leaf_47_wb_clk_i _03115_ _01418_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12458__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14767_ net1186 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XANTENNA__08638__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ net2527 net222 net469 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16506_ clknet_leaf_102_wb_clk_i net3009 _00369_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_13718_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] _04027_ vssd1 vssd1 vccd1 vccd1
+ _04038_ sky130_fd_sc_hd__nand2_1
XANTENNA__11642__A1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10445__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17486_ clknet_leaf_53_wb_clk_i _03046_ _01349_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14698_ net1406 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16437_ clknet_leaf_77_wb_clk_i _02065_ _00300_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_13649_ _03806_ _03969_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13395__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16368_ clknet_leaf_66_wb_clk_i net1776 _00236_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09994__C net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18107_ net1481 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_82_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15319_ net1244 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XANTENNA__12193__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16299_ clknet_leaf_111_wb_clk_i _01933_ _00167_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09068__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18038_ net1428 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_2_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout317 _07975_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_2
X_09811_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[7\] net862 vssd1
+ vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and3_1
Xfanout328 _03750_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
Xfanout339 _06982_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17873__CLK clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08700__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09742_ net1007 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[10\] net864
+ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18156__1530 vssd1 vssd1 vccd1 vccd1 _18156__1530/HI net1530 sky130_fd_sc_hd__conb_1
X_09673_ net1091 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[11\] net869
+ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__and3_1
XANTENNA__09234__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13870__A2 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_A _07948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17103__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[29\] net663 net632 team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09531__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\] net746 net745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a22o_1
XANTENNA__08629__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12368__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A _08021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10436__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08486_ net1112 net1115 net1107 net1109 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__and4b_4
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13386__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112__1486 vssd1 vssd1 vccd1 vccd1 _18112__1486/HI net1486 sky130_fd_sc_hd__conb_1
X_09107_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] net726 net687 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[17\]
+ _05352_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09038_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[18\] net716 net697 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[18\]
+ _05284_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold360 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12831__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12897__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[9\] vssd1 vssd1 vccd1 vccd1
+ net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[6\] vssd1 vssd1 vccd1 vccd1
+ net2009 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net323 _07247_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09706__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout840 team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1
+ net840 sky130_fd_sc_hd__clkbuf_4
Xfanout851 net854 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
Xfanout862 _04754_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_4
Xfanout873 net874 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
Xfanout884 _04744_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout895 _04738_ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__buf_4
X_12951_ team_01_WB.instance_to_wrap.a1.ADR_I\[10\] net606 net588 _03640_ vssd1 vssd1
+ vccd1 vccd1 _02218_ sky130_fd_sc_hd__a22o_1
Xhold1060 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 _03417_ vssd1 vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net3183 net191 net475 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__mux2_1
Xhold1082 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
X_15670_ net1260 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
X_12882_ net2886 net607 net589 _03590_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
Xhold1093 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08983__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14621_ net1369 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ net679 _07344_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__nand2_1
XANTENNA__12278__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17340_ clknet_leaf_20_wb_clk_i _02900_ _01203_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14552_ net1334 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XANTENNA__10427__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11764_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[24\] _07861_ vssd1 vssd1
+ vccd1 vccd1 _07898_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ _03852_ _03854_ _03855_ _03769_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10715_ _06866_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__nor2_1
XANTENNA__13898__A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17271_ clknet_leaf_9_wb_clk_i _02831_ _01134_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14483_ net1400 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
X_11695_ team_01_WB.instance_to_wrap.cpu.K0.count\[1\] team_01_WB.instance_to_wrap.cpu.K0.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11910__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ clknet_leaf_42_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[3\]
+ _00090_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17746__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13377__B2 team_01_WB.instance_to_wrap.cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13434_ _03781_ _03786_ _03780_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10646_ _05620_ _05583_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16153_ net1332 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ net486 _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ _04959_ _06838_ _06840_ _06839_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08504__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ net1273 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net2806 net216 net427 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux2_1
X_16084_ net1403 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__inv_2
X_13296_ net1756 net808 net803 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[28\] vssd1
+ vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17896__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15035_ net1298 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12247_ net2997 net255 net437 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__mux2_1
XANTENNA__12741__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12178_ net2091 net222 net445 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11560__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17126__CLK clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _06996_ _07294_ _07295_ net330 vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16986_ clknet_leaf_34_wb_clk_i _02546_ _00849_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09054__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15937_ net1340 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__inv_2
XANTENNA__08859__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15868_ net1396 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__inv_2
XANTENNA__09989__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17607_ clknet_leaf_130_wb_clk_i _03167_ _01470_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14819_ net1353 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XANTENNA__13065__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12188__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15799_ net1239 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10418__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ net2918 net3081 net1038 vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
X_17538_ clknet_leaf_0_wb_clk_i _03098_ _01401_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11615__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08271_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[85\] team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[77\]
+ net1045 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17469_ clknet_leaf_14_wb_clk_i _03029_ _01332_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09036__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08414__B _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14317__B1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09229__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18054__1616 vssd1 vssd1 vccd1 vccd1 net1616 _18054__1616/LO sky130_fd_sc_hd__conb_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12651__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09526__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08430__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\] net721 net718 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[10\]
+ _05980_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a221o_1
XANTENNA__17619__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1398_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[11\] net733 _05917_ _05918_
+ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08607_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[29\] net726 _04856_
+ _04859_ _04860_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12098__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13056__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09587_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] net709 net757 vssd1
+ vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout823_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17769__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ net975 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\] net936 vssd1
+ vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and3_1
XANTENNA__10200__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12826__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ net1108 net1115 net1112 net1106 vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_46_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13359__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[25\] net651 _04765_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[25\] _06763_ vssd1 vssd1 vccd1
+ vccd1 _06764_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11480_ _07729_ _07732_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire559 _05618_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_4
XFILLER_0_85_1642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10431_ _06684_ _06689_ _06693_ _06694_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__or4_4
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13150_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[84\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[92\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10362_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\] net693 net686 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__a22o_1
XANTENNA__09139__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ net494 _08011_ _08017_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__and3_4
XFILLER_0_108_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17149__CLK clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11966__A team_01_WB.instance_to_wrap.cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[0\] net623 _06554_ _06555_
+ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a2111o_1
X_13081_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[13\] net1030 vssd1 vssd1 vccd1
+ vccd1 _03708_ sky130_fd_sc_hd__or2_1
XANTENNA__14342__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[16\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ net1985 net292 net464 vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XANTENNA__09436__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[27\] vssd1 vssd1 vccd1 vccd1
+ net1806 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12885__A3 _03592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ clknet_leaf_45_wb_clk_i _02400_ _00703_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16173__CLK clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17299__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout670 _04729_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_8
Xfanout681 _04717_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_4
Xfanout692 net694 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_4
X_16771_ clknet_leaf_119_wb_clk_i _02331_ _00634_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13983_ _03556_ _04169_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__nor2_1
XANTENNA__11905__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15722_ net1198 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12934_ net1026 _07535_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15653_ net1232 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13047__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12865_ net1034 _03575_ _03576_ net1161 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a211o_1
XANTENNA__09602__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14604_ net1399 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
X_11816_ net679 _07223_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15584_ net1269 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12796_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[31\] _07869_ net373 vssd1
+ vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17323_ clknet_leaf_61_wb_clk_i _02883_ _01186_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14535_ net1320 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11747_ net3050 net238 net479 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11640__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17254_ clknet_leaf_140_wb_clk_i _02814_ _01117_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14466_ net1390 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11678_ net1636 net1160 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16205_ clknet_4_8__leaf_wb_clk_i _01872_ _00073_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13417_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[27\] team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\]
+ net591 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10629_ _06277_ net544 vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17185_ clknet_leaf_138_wb_clk_i _02745_ _01048_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14397_ net1329 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16136_ net1321 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__inv_2
X_13348_ net8 net798 net593 net3030 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09049__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13567__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16067_ net1401 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__inv_2
XANTENNA__15348__A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12471__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__A_N _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ net1788 net810 net597 team_01_WB.instance_to_wrap.a1.ADR_I\[12\] vssd1 vssd1
+ vccd1 vccd1 _01995_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09726__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13522__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ net1223 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__16516__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14078__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16969_ clknet_leaf_49_wb_clk_i _02529_ _00832_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09510_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[9\] net735 net685 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a22o_1
XANTENNA__16666__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18111__1485 vssd1 vssd1 vccd1 vccd1 _18111__1485/HI net1485 sky130_fd_sc_hd__conb_1
X_09441_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\] net742 net741 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a22o_1
XANTENNA__13038__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13589__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10020__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09372_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[13\] net741 _05623_ _05627_
+ _05632_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14250__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ net3212 net3178 net1049 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12646__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A _07893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13331__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08254_ net3002 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[94\] net1039 vssd1 vssd1
+ vccd1 vccd1 _03493_ sky130_fd_sc_hd__mux2_1
XANTENNA__09009__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08425__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08185_ _04564_ _04572_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout404_A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13761__A1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11772__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10690__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1313_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13277__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09708_ net981 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[10\] net928 vssd1
+ vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17591__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ _05485_ _06606_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nor2_1
XANTENNA__09350__D1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13029__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ net1135 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[11\] net954
+ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15721__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12650_ net2633 net273 net391 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09248__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14241__A2 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11601_ net496 _07815_ net2255 net838 vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12581_ net2212 net216 net399 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__mux2_1
XANTENNA__12556__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ net2803 _04455_ _04457_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ team_01_WB.instance_to_wrap.cpu.f0.i\[14\] _07707_ vssd1 vssd1 vccd1 vccd1
+ _07768_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[78\] _04229_ _04247_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[86\]
+ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__a22o_1
X_11463_ _04469_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ net2240 net2125 net818 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
X_10414_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[26\] net935
+ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and3_1
XANTENNA__11212__C1 _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18135__1509 vssd1 vssd1 vccd1 vccd1 _18135__1509/HI net1509 sky130_fd_sc_hd__conb_1
X_14182_ net793 _04233_ _04249_ _04279_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__or4_1
X_11394_ _07288_ _07551_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__nor3_1
XFILLER_0_123_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15168__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[101\] team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ net822 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
X_10345_ _05278_ _05347_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12291__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09166__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[18\] _03695_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__mux2_1
X_17941_ clknet_leaf_106_wb_clk_i _03491_ _01761_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[100\]
+ sky130_fd_sc_hd__dfstp_1
X_10276_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[0\] net888 vssd1
+ vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__and3_1
XANTENNA__08070__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09184__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ net3225 net256 net464 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
Xfanout1410 net1411 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__buf_4
XFILLER_0_104_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17872_ clknet_leaf_100_wb_clk_i _03422_ _01692_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14800__A net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17934__CLK clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16823_ clknet_leaf_24_wb_clk_i _02383_ _00686_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13268__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16754_ clknet_leaf_40_wb_clk_i _02314_ _00617_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13966_ team_01_WB.instance_to_wrap.cpu.LCD0.currentState\[0\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ net584 vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12917_ net1031 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[19\] vssd1 vssd1 vccd1
+ vccd1 _03616_ sky130_fd_sc_hd__or2_1
X_15705_ net1237 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
X_16685_ clknet_leaf_55_wb_clk_i _02245_ _00548_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09332__C net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ net2935 net796 vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[10\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053__1615 vssd1 vssd1 vccd1 vccd1 net1615 _18053__1615/LO sky130_fd_sc_hd__conb_1
XFILLER_0_5_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15631__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15636_ net1241 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
X_12848_ net2199 net273 net367 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12974__B net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14232__A2 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08447__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12466__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15567_ net1201 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
X_12779_ net1800 net218 net375 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ net1396 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
X_17306_ clknet_leaf_36_wb_clk_i _02866_ _01169_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15498_ net1202 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14449_ net1392 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17237_ clknet_leaf_9_wb_clk_i _02797_ _01100_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10006__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13743__A1 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09947__B1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold904 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ clknet_leaf_25_wb_clk_i _02728_ _01031_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17464__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold915 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[105\] vssd1 vssd1 vccd1 vccd1
+ net2542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16119_ net1369 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__inv_2
Xhold937 _03413_ vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold948 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09990_ net1138 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\] net954 vssd1
+ vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__and3_1
X_17099_ clknet_leaf_60_wb_clk_i _02659_ _00962_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold959 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[87\] vssd1 vssd1 vccd1 vccd1
+ net2575 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08941_ _05166_ _05201_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ _05099_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1604 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1626 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3242 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1637 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net3253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1648 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net3264
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout187_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11809__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08686__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout354_A net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1096_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15541__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ net548 _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13026__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14223__A2 _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08438__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ net1155 net576 net577 net582 vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10685__A _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12376__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout619_A _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1263_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10245__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ net2867 net2747 net1052 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09286_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[15\] net576 _05242_ vssd1 vssd1
+ vccd1 vccd1 _05550_ sky130_fd_sc_hd__a21o_1
XANTENNA__09650__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17807__CLK clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ net2330 net2205 net1044 vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08168_ _04563_ team_01_WB.instance_to_wrap.cpu.K0.code\[3\] team_01_WB.instance_to_wrap.cpu.K0.code\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__or3b_2
XFILLER_0_107_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_108_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout988_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08610__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ _04465_ team_01_WB.instance_to_wrap.cpu.f0.num\[24\] team_01_WB.instance_to_wrap.cpu.f0.num\[15\]
+ _04472_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13000__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17957__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10130_ net986 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[2\] _04666_ vssd1
+ vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10061_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[3\] net919 vssd1
+ vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__and3_1
XANTENNA__09714__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13820_ team_01_WB.instance_to_wrap.cpu.c0.count\[6\] _04112_ vssd1 vssd1 vccd1 vccd1
+ _04113_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ net1666 _04063_ net783 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08677__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _06922_ _06926_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13670__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10298__C net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12702_ net2494 net235 net383 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
X_16470_ clknet_leaf_85_wb_clk_i _02098_ _00333_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_13682_ _03784_ _03785_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _05138_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15421_ net1277 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12633_ net2982 net209 net393 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12286__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10595__A team_01_WB.instance_to_wrap.cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18140_ net1514 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
XFILLER_0_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15352_ net1242 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
X_12564_ _08008_ _08012_ net488 vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__and3_4
XFILLER_0_4_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10787__A1 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14303_ team_01_WB.instance_to_wrap.cpu.LCD0.cnt_20ms\[9\] _04445_ net1366 vssd1
+ vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11515_ _07754_ _07756_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18071_ net1445 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15283_ net1177 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
X_12495_ net1891 net294 net414 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17022_ clknet_leaf_2_wb_clk_i _02582_ _00885_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13725__A1 _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14234_ _04384_ _04386_ _04388_ _04390_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__or4_1
X_11446_ net486 _07698_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__nand2b_1
X_18110__1484 vssd1 vssd1 vccd1 vccd1 _18110__1484/HI net1484 sky130_fd_sc_hd__conb_1
XFILLER_0_85_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14165_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[74\] _04229_ _04242_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[2\]
+ _04313_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a221o_1
XANTENNA__11200__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11377_ _06778_ _07123_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08512__B net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[118\] net1904 net819 vssd1 vssd1
+ vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
X_10328_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__inv_2
X_14096_ net792 net791 _04237_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__and3_4
XANTENNA__09327__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\] net836 net356 _03684_ vssd1
+ vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a22o_1
X_17924_ clknet_leaf_82_wb_clk_i _03474_ _01744_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ net579 _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1240 net1245 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
Xfanout1251 net1253 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17855_ clknet_leaf_102_wb_clk_i _03405_ _01675_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1262 net1264 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
Xfanout1273 net1276 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1284 net1285 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_2
Xfanout1295 net1296 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__clkbuf_4
X_16806_ clknet_leaf_141_wb_clk_i _02366_ _00669_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_17786_ clknet_leaf_114_wb_clk_i _03344_ _01607_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14998_ net1258 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XANTENNA__09062__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13661__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16737_ clknet_leaf_138_wb_clk_i _02297_ _00600_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08668__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13949_ net1163 net1057 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[30\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[30\] sky130_fd_sc_hd__and3b_1
XFILLER_0_18_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16668_ clknet_leaf_115_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[22\]
+ _00531_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09997__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14205__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12196__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15619_ net1219 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16599_ clknet_leaf_58_wb_clk_i _02227_ _00462_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09140_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[17\] net608 _05382_
+ _05389_ _05396_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11424__C1 _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09071_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[18\] net638 _05312_ _05313_
+ _05316_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08703__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold701 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold712 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold723 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold734 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10671__C _06933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold767 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[15\] vssd1 vssd1 vccd1 vccd1
+ net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[5\] net645 _06224_ _06226_
+ _06229_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a2111o_1
Xhold789 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__A1 _06992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08924_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[21\] net665 net653 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a22o_1
XANTENNA__15536__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1401 team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net3017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12879__B _07600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_141_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1412 team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3028 sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[20\] net882 vssd1
+ vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__and3_1
Xhold1423 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout471_A _08010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1434 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net3050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\] vssd1 vssd1 vccd1 vccd1
+ net3061 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1456 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net3072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1467 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net3083 sky130_fd_sc_hd__dlygate4sd3_1
X_08786_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[22\] net644 net622 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a22o_1
Xhold1478 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[81\] vssd1 vssd1 vccd1 vccd1
+ net3094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1489 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net3105 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13652__A0 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08659__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18134__1508 vssd1 vssd1 vccd1 vccd1 _18134__1508/HI net1508 sky130_fd_sc_hd__conb_1
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1380_A net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09871__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ net1069 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[13\] net850
+ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09700__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09338_ net1081 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[14\] net892
+ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12834__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ net1071 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[15\] net891
+ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13707__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ _05963_ _06029_ _07498_ net345 vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12280_ net2257 net255 net432 vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__mux2_1
XANTENNA__09709__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10862__B _06933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09387__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ _06869_ _07481_ _07482_ _07494_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__a31o_2
XFILLER_0_82_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11162_ _07422_ _07423_ _07425_ _07421_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__a211o_2
X_18052__1614 vssd1 vssd1 vccd1 vccd1 net1614 _18052__1614/LO sky130_fd_sc_hd__conb_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ _06373_ _06374_ _06375_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15446__A net1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15970_ net1332 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__inv_2
XANTENNA__14350__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _05852_ _06071_ net504 vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08986__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[4\] net663 _06282_ _06285_
+ _06294_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a2111o_1
X_14921_ net1214 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08898__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[23\] vssd1 vssd1 vccd1 vccd1
+ net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 team_01_WB.instance_to_wrap.cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1
+ net1677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17640_ clknet_leaf_45_wb_clk_i _03200_ _01503_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold72 team_01_WB.instance_to_wrap.cpu.f0.write_data\[14\] vssd1 vssd1 vccd1 vccd1
+ net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 _01959_ vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1350 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
Xhold94 net146 vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16727__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ net563 _07772_ _04103_ net786 vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a31o_1
X_14783_ net1407 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
X_17571_ clknet_leaf_133_wb_clk_i _03131_ _01434_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11995_ net2472 net261 net469 vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
XANTENNA_output119_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11913__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15181__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13734_ net563 _04019_ _04049_ _04050_ net786 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a311o_1
XFILLER_0_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16522_ clknet_leaf_81_wb_clk_i _02150_ _00385_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10946_ _07162_ _07167_ net509 vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09862__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16453_ clknet_leaf_80_wb_clk_i net1658 _00316_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_13665_ net769 _03991_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09610__C net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _07004_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__nand2_1
XANTENNA__16877__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10209__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08507__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12616_ net2549 net248 net395 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
X_15404_ net1263 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
X_16384_ clknet_leaf_83_wb_clk_i _00001_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ net966 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\] _03934_ _03935_
+ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
XANTENNA__09614__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18123_ net1497 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
X_15335_ net1180 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
X_12547_ net2444 net278 net404 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08822__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12744__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18054_ net1616 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
X_15266_ net1266 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
X_12478_ net2145 net219 net411 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[125\] _04233_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[109\]
+ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__a22o_1
X_17005_ clknet_leaf_19_wb_clk_i _02565_ _00868_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11429_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[7\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[6\]
+ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[5\] team_01_WB.instance_to_wrap.cpu.DM0.data_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15197_ net1282 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11185__A1 _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ net1892 net585 _04308_ net1170 vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09057__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10393__C1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16257__CLK clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15356__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[3\] team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__and2_2
XFILLER_0_20_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17502__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17907_ clknet_leaf_81_wb_clk_i _03457_ _01727_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11488__A2 _07734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_2
Xfanout1081 net1088 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_2
X_08640_ net583 _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__or2_1
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_2
X_17838_ clknet_leaf_91_wb_clk_i _03389_ _01659_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12437__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[30\] net652 net629 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[30\]
+ _04834_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a221o_1
XANTENNA__17652__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__A0 _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17769_ clknet_leaf_97_wb_clk_i _03327_ _01590_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10448__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08417__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09123_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[17\] net852 vssd1
+ vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__and3_1
XANTENNA__12654__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout317_A _07975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1059_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ net1004 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[18\] net842 vssd1
+ vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09529__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17032__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold520 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[29\] vssd1 vssd1 vccd1 vccd1
+ net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1 vccd1 net2158
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold553 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold564 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold575 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[72\] vssd1 vssd1 vccd1 vccd1
+ net2202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold597 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11794__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[5\] net858 vssd1
+ vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08907_ net1074 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[21\] net858
+ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__and3_1
XANTENNA__12676__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ net1018 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[6\] net888 vssd1
+ vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout853_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 team_01_WB.instance_to_wrap.cpu.f0.num\[6\] vssd1 vssd1 vccd1 vccd1 net2858
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[20\] net856
+ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__and3_1
XANTENNA__10203__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1253 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[70\] vssd1 vssd1 vccd1 vccd1
+ net2869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1264 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 _02071_ vssd1 vssd1 vccd1 vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1286 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1297 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08769_ _05030_ _05031_ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__or3_1
XANTENNA__12829__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10439__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ net509 _07063_ net520 vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11780_ net2672 net229 net479 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11100__A1 _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09844__A2 _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10731_ _06952_ _06978_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__nor2_2
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09430__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ _03799_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10662_ _05419_ _06925_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ net1919 net192 net419 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ team_01_WB.instance_to_wrap.cpu.f0.num\[17\] net329 net353 net1894 vssd1
+ vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10593_ _04725_ _06847_ _06850_ net1155 vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__a22o_1
XANTENNA__14345__A team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[13\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ net1250 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
X_12332_ _07834_ _07843_ _07840_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[11\] vssd1
+ vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_134_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15051_ net1204 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_12263_ net2522 net296 net438 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14002_ _04170_ _04177_ _04179_ _04186_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o31a_1
XFILLER_0_82_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11214_ _07464_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12194_ net2648 net261 net445 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11908__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _07406_ _07408_ net541 vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__mux2_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10390__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_37_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17675__CLK clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15953_ net1330 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__inv_2
X_11076_ net541 _07339_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__nor2_1
XANTENNA__09605__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net1022 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[4\] net894 vssd1
+ vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and3_1
X_14904_ net1306 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
X_15884_ net1352 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__inv_2
XANTENNA__10142__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17623_ clknet_leaf_11_wb_clk_i _03183_ _01486_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14835_ net1339 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XANTENNA__12739__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13616__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13424__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17554_ clknet_leaf_23_wb_clk_i _03114_ _01417_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08099__B2 _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__A1 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14766_ net1184 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
X_11978_ net2733 net228 net467 vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09835__A2 _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16505_ clknet_leaf_99_wb_clk_i _02133_ _00368_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[117\]
+ sky130_fd_sc_hd__dfstp_1
X_13717_ _04022_ _04036_ _04558_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__a21oi_1
X_10929_ _07144_ _07179_ _07189_ _06970_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__a22o_1
XANTENNA__09340__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14697_ net1402 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
X_17485_ clknet_leaf_21_wb_clk_i _03045_ _01348_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18205__1579 vssd1 vssd1 vccd1 vccd1 _18205__1579/HI net1579 sky130_fd_sc_hd__conb_1
XANTENNA__10850__A0 _05515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16436_ clknet_leaf_103_wb_clk_i _02064_ _00299_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13648_ net968 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] _03978_ _03979_
+ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16367_ clknet_leaf_66_wb_clk_i net1838 _00235_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12474__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13579_ net186 _07917_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18106_ net1480 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
X_15318_ net1260 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16298_ clknet_leaf_109_wb_clk_i _01932_ _00166_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18037_ net1427 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_2_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15249_ net1195 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap916_A _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18133__1507 vssd1 vssd1 vccd1 vccd1 _18133__1507/HI net1507 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout307 net310 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
X_09810_ net1097 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[7\] net898 vssd1
+ vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__and3_1
XANTENNA__08574__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout329 _03750_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10381__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ net1086 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[10\] net857
+ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09672_ net1090 team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[11\] net858
+ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10023__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10133__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[29\] net637 _04765_
+ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[29\] _04885_ vssd1 vssd1 vccd1
+ vccd1 _04887_ sky130_fd_sc_hd__a221o_1
XANTENNA__09812__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13607__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12649__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10958__A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08554_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[30\] net724 net684 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a22o_1
XANTENNA__09287__A0 _05549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13083__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13946__A_N net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08428__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08485_ net1003 net872 vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__and2_4
X_18051__1613 vssd1 vssd1 vccd1 vccd1 net1613 _18051__1613/LO sky130_fd_sc_hd__conb_1
XANTENNA__11633__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_A _08023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1176_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09039__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12384__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17548__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _05365_ _05366_ _05367_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09259__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _05297_ _05298_ _05299_ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13543__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16572__CLK clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__S net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__A1 team_01_WB.instance_to_wrap.cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold394 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[5\] vssd1 vssd1 vccd1 vccd1
+ net2010 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout830 net832 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10372__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout841 team_01_WB.instance_to_wrap.cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1
+ net841 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout852 net855 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_4
X_09939_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[23\]\[5\] net686 _06200_ _06201_
+ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__a2111o_1
Xfanout863 net866 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_4
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
XANTENNA__11029__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout885 net889 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_4
X_12950_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[10\] net1055 net365 _03639_
+ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a22o_1
Xfanout896 net900 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_4
XANTENNA__15724__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11321__B2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1061 team_01_WB.instance_to_wrap.cpu.f0.num\[26\] vssd1 vssd1 vccd1 vccd1 net2677
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net2895 net194 net477 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__mux2_1
Xhold1072 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ net366 _03588_ _03589_ net1056 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a32o_1
Xhold1083 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\] vssd1 vssd1 vccd1 vccd1
+ net2699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12559__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1094 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[15\] vssd1 vssd1 vccd1 vccd1
+ net2710 sky130_fd_sc_hd__dlygate4sd3_1
X_11832_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[12\] _07853_ vssd1 vssd1
+ vccd1 vccd1 _07954_ sky130_fd_sc_hd__xnor2_1
X_14620_ net1385 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14271__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ net1335 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09160__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ net2893 net232 net481 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[22\] _05064_ _03843_ _03842_
+ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a31oi_1
X_10714_ _06856_ _06858_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_49_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17270_ clknet_leaf_30_wb_clk_i _02830_ _01133_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14482_ net1380 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
XANTENNA__13898__B net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11694_ net3107 net154 team_01_WB.instance_to_wrap.cpu.K0.next_state vssd1 vssd1
+ vccd1 vccd1 _03258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16221_ clknet_leaf_43_wb_clk_i team_01_WB.instance_to_wrap.cpu.c0.next_count\[2\]
+ _00089_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.c0.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_13433_ _03784_ _03785_ _03783_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a21o_1
XANTENNA__12294__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645_ _05551_ _05515_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16152_ net1323 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13364_ _04503_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _07680_ vssd1 vssd1
+ vccd1 vccd1 _03749_ sky130_fd_sc_hd__a21oi_1
X_10576_ _04906_ _04907_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__nor2_2
XFILLER_0_10_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap1169 _07837_ vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_2
X_15103_ net1294 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
X_12315_ net1852 net280 net427 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
X_16083_ net1400 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__inv_2
X_13295_ net1816 net808 net803 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[29\] vssd1
+ vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15034_ net1305 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
X_12246_ net2843 net220 net437 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_91_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11638__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12177_ net2082 net229 net443 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11560__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11128_ _07106_ _07391_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nand2_1
XANTENNA__09335__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16985_ clknet_leaf_14_wb_clk_i _02545_ _00848_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15936_ net1340 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__inv_2
X_11059_ _07004_ _07321_ _07322_ _07079_ _07319_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__a221o_1
XANTENNA__10115__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12977__B _07456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09632__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15867_ net1393 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12469__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17606_ clknet_leaf_141_wb_clk_i _03166_ _01469_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14818_ net1354 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15798_ net1304 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__inv_2
XANTENNA__14262__B1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17537_ clknet_leaf_137_wb_clk_i _03097_ _01400_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14749_ net1311 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10823__A0 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08270_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[86\] net2600 net1040 vssd1 vssd1
+ vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17468_ clknet_leaf_13_wb_clk_i _03028_ _01331_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16419_ clknet_leaf_100_wb_clk_i _02047_ _00282_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17399_ clknet_leaf_11_wb_clk_i _02959_ _01262_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09441__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10051__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11551__B2 _07731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout384_A _03568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\] net700 _05986_ _05987_
+ net712 vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10106__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__B _07585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09542__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17220__CLK clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[11\] net751 net704 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a22o_1
XANTENNA__12379__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1293_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_A _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[29\] net744 _04855_ _04863_
+ _04864_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _05839_ _05844_ _05848_ _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__or4_4
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14253__B1 _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ net1124 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[30\] net953
+ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__and3_1
XANTENNA__11067__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout816_A _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08468_ net1086 net907 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__and2_2
XFILLER_0_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13359__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08399_ net1147 net1149 net1151 net1153 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_11_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13003__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10430_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\] net745 net738 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[26\]
+ _06680_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08786__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10361_ net985 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[27\] net938 vssd1
+ vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12842__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12100_ team_01_WB.instance_to_wrap.cpu.IG0.Instr\[10\] team_01_WB.instance_to_wrap.cpu.IG0.Instr\[9\]
+ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__and2b_2
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ _05685_ _07807_ _03704_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11966__B team_01_WB.instance_to_wrap.cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10292_ net1020 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[0\] net899 vssd1
+ vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__and3_1
X_12031_ net2728 net295 net466 vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold180 _01973_ vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 team_01_WB.instance_to_wrap.cpu.f0.write_data\[19\] vssd1 vssd1 vccd1 vccd1
+ net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18204__1578 vssd1 vssd1 vccd1 vccd1 _18204__1578/HI net1578 sky130_fd_sc_hd__conb_1
XFILLER_0_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout660 net661 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13673__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout671 _04729_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16770_ clknet_leaf_144_wb_clk_i _02330_ _00633_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13982_ _04167_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__nor2_1
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_6
XANTENNA__08994__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15721_ net1214 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
X_12933_ net1849 net605 net587 _03627_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a22o_1
XANTENNA__12289__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08710__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13047__A1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15652_ net1269 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
X_12864_ net1034 team_01_WB.instance_to_wrap.cpu.f0.write_i vssd1 vssd1 vccd1 vccd1
+ _03576_ sky130_fd_sc_hd__nor2_1
XANTENNA__14244__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18132__1506 vssd1 vssd1 vccd1 vccd1 _18132__1506/HI net1506 sky130_fd_sc_hd__conb_1
X_14603_ net1371 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
X_11815_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[15\] _07855_ vssd1 vssd1
+ vccd1 vccd1 _07940_ sky130_fd_sc_hd__xnor2_1
X_15583_ net1295 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
XANTENNA_output101_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12795_ _07842_ _07845_ net489 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and3_4
XANTENNA__11921__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17322_ clknet_leaf_43_wb_clk_i _02882_ _01185_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14534_ net1331 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
X_11746_ net781 _07881_ _07882_ _07883_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__a22o_2
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17863__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17253_ clknet_leaf_133_wb_clk_i _02813_ _01116_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14465_ net1390 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
X_11677_ net1719 net1160 vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16204_ clknet_leaf_105_wb_clk_i _01871_ _00072_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10628_ _06245_ _06211_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__nand2b_1
X_13416_ _03767_ _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14396_ net1329 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
X_17184_ clknet_leaf_140_wb_clk_i _02744_ _01047_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16135_ net1330 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__inv_2
X_13347_ net9 net799 net594 net2994 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13770__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12752__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10559_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[8\]\[24\] net648 net612 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13278_ net79 net810 net597 net1913 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
X_16066_ net1405 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08529__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net2250 net309 net442 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
X_15017_ net1205 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
X_18050__1612 vssd1 vssd1 vccd1 vccd1 net1612 _18050__1612/LO sky130_fd_sc_hd__conb_1
XANTENNA__11533__A1 team_01_WB.instance_to_wrap.cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17243__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09065__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16968_ clknet_leaf_45_wb_clk_i _02528_ _00831_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09362__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ net1353 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__inv_2
XANTENNA__12199__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16899_ clknet_leaf_120_wb_clk_i _02459_ _00762_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17393__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[12\] net706 _05691_
+ _05692_ _05702_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10301__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11049__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08409__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13589__A2 _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09371_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[13\] net730 net702 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08322_ net2695 net2686 net1047 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_89_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08706__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13331__B net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ net3076 net2829 net1045 vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ _04553_ _04571_ _04575_ _04564_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11874__A1_N net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08768__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12662__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14443__A net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1139_A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09537__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10690__B _06953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A _03742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11889__A1_N team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1306_A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1414_A team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ net1132 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[10\] net943
+ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__and3_1
XANTENNA__09703__C net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09638_ net1137 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[11\] net952
+ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__and3_1
XANTENNA__14226__B1 _04281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16760__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ net1129 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[8\] net948 vssd1
+ vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12837__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ team_01_WB.instance_to_wrap.cpu.DM0.data_i\[26\] net572 vssd1 vssd1 vccd1
+ vccd1 _07815_ sky130_fd_sc_hd__nand2_1
XANTENNA__11741__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12580_ net2614 net278 net400 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09653__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11531_ team_01_WB.instance_to_wrap.cpu.f0.i\[15\] _07766_ _07767_ _07731_ vssd1
+ vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14250_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[46\] _04268_ _04281_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[30\]
+ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a221o_1
X_11462_ team_01_WB.instance_to_wrap.cpu.f0.i\[18\] _07713_ vssd1 vssd1 vccd1 vccd1
+ _07715_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[33\] net3089 net829 vssd1 vssd1
+ vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
XANTENNA__13668__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ net1117 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[26\] net948
+ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ _04225_ net790 net788 _04261_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a31o_1
XANTENNA__12572__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11393_ _07324_ _07535_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12960__B1 team_01_WB.instance_to_wrap.cpu.RU0.state\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13132_ net2524 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[110\] net819 vssd1 vssd1
+ vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XANTENNA_input62_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08989__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17266__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10344_ _05417_ _05483_ _05418_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11188__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17940_ clknet_leaf_81_wb_clk_i net2483 _01760_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_13063_ _05344_ net570 net358 vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10275_ net1102 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[0\] net849 vssd1
+ vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10318__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12014_ net3047 net221 net464 vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
Xfanout1400 net1413 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__buf_4
Xfanout1411 net1412 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__buf_4
X_17871_ clknet_leaf_102_wb_clk_i _03421_ _01691_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11916__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16822_ clknet_leaf_29_wb_clk_i _02382_ _00685_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 _08025_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09182__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16753_ clknet_leaf_24_wb_clk_i _02313_ _00616_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ net584 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__inv_2
XANTENNA__09613__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15704_ net1254 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
X_12916_ net1027 _07625_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16684_ clknet_leaf_61_wb_clk_i _02244_ _00547_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10121__A _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14217__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[9\] net797 vssd1 vssd1 vccd1 vccd1
+ team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedInstr\[9\] sky130_fd_sc_hd__and2_1
X_15635_ net1187 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XANTENNA__12747__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ net2166 net248 net368 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13432__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ net1230 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09644__B1 _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12778_ net3022 net280 net376 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17305_ clknet_leaf_125_wb_clk_i _02865_ _01168_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14517_ net1409 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ net2512 net197 net481 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15497_ net1215 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17236_ clknet_leaf_7_wb_clk_i _02796_ _01099_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14448_ net1390 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11887__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11203__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12482__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17167_ clknet_leaf_93_wb_clk_i _02727_ _01030_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14379_ net1328 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold905 team_01_WB.instance_to_wrap.cpu.RU0.state\[2\] vssd1 vssd1 vccd1 vccd1 net2521
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10557__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold916 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _02129_ vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09357__A _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16118_ net1359 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
X_17098_ clknet_leaf_42_wb_clk_i _02658_ _00961_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold949 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10962__C1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11098__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ _05166_ _05202_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16049_ net1364 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__inv_2
XANTENNA__16633__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17759__CLK clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09175__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_131_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08871_ _05133_ _05134_ net578 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__mux2_1
XANTENNA__10015__B _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1605 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net3221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1616 team_01_WB.instance_to_wrap.cpu.RF0.registers\[13\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net3232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1627 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net3243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1638 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net3254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1649 team_01_WB.instance_to_wrap.cpu.c0.count\[13\] vssd1 vssd1 vccd1 vccd1 net3265
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16783__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10031__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14208__B1 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09423_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__inv_2
XANTENNA__09820__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__A2_N net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17139__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[14\] net669 _05613_ _05617_
+ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_34_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1089_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13431__A1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10685__B _06867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08305_ net3111 net3079 net1051 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[15\] net666 _05545_ _05548_
+ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o22a_4
X_18203__1577 vssd1 vssd1 vccd1 vccd1 _18203__1577/HI net1577 sky130_fd_sc_hd__conb_1
XANTENNA_fanout514_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1256_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[120\] net1680 net1039 vssd1 vssd1
+ vccd1 vccd1 _03511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16163__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ net1755 net553 _04569_ net1065 vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__a22o_1
XANTENNA__12392__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10548__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ _04488_ team_01_WB.instance_to_wrap.cpu.f0.i\[29\] _04461_ team_01_WB.instance_to_wrap.cpu.f0.num\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_105_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout883_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08602__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18131__1505 vssd1 vssd1 vccd1 vccd1 _18131__1505/HI net1505 sky130_fd_sc_hd__conb_1
XFILLER_0_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10060_ net1145 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[3\] net952 vssd1
+ vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09433__C net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ net485 _07719_ _04060_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__a31o_1
X_10962_ _05348_ _07224_ _07225_ net346 vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13670__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12701_ net2722 net202 net385 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13681_ _04005_ _04004_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] net968
+ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12567__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ _06878_ _06919_ _06921_ _06928_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__a31o_1
X_15420_ net1277 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ net2682 net193 net391 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16506__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ net3099 net213 net406 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15351_ net1238 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11514_ _07716_ _07724_ _07734_ team_01_WB.instance_to_wrap.cpu.f0.i\[20\] vssd1
+ vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__a31o_1
X_14302_ _04445_ _04446_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18070_ net1444 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
X_12494_ net2794 net308 net414 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__mux2_1
X_15282_ net1174 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
X_17021_ clknet_leaf_127_wb_clk_i _02581_ _00884_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11445_ _07682_ team_01_WB.instance_to_wrap.cpu.f0.state\[6\] _04619_ vssd1 vssd1
+ vccd1 vccd1 _07698_ sky130_fd_sc_hd__or3b_1
XFILLER_0_62_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14233_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[5\] _04242_ _04267_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[13\]
+ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16656__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10539__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__A team_01_WB.instance_to_wrap.cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17901__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _04320_ _04321_ _04322_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11376_ net344 _07626_ _07628_ _07639_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09608__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10327_ net554 _06590_ team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\] net760
+ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a2bb2o_1
X_13115_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[119\] net2034 net824 vssd1 vssd1
+ vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14095_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[48\] _04255_ _04256_ team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[104\]
+ _04254_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13046_ team_01_WB.instance_to_wrap.cpu.f0.write_data\[24\] _03683_ net1030 vssd1
+ vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__mux2_1
X_17923_ clknet_leaf_82_wb_clk_i _03473_ _01743_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14150__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ net579 _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1230 net1235 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13427__A team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1241 net1245 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_4
X_17854_ clknet_leaf_98_wb_clk_i _03404_ _01674_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_10189_ _06414_ net530 vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__and2_1
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_4
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_4
Xfanout1274 net1276 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_4
Xfanout1285 net1301 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16805_ clknet_leaf_129_wb_clk_i _02365_ _00668_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1296 net1301 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_2
XANTENNA__09343__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17785_ clknet_leaf_113_wb_clk_i _03343_ _01606_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14997_ net1177 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XANTENNA__10489__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15642__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16736_ clknet_leaf_142_wb_clk_i _02296_ _00599_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ net1164 net1057 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[29\] vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[29\] sky130_fd_sc_hd__and3b_1
XFILLER_0_57_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09640__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16667_ clknet_leaf_106_wb_clk_i team_01_WB.instance_to_wrap.cpu.RU0.next_FetchedData\[21\]
+ _00530_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.data_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11672__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ team_01_WB.instance_to_wrap.cpu.RU0.state\[6\] net1059 net1165 vssd1 vssd1
+ vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RU0.next_dhit sky130_fd_sc_hd__o21ba_1
XFILLER_0_9_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15618_ net1289 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16186__CLK clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16598_ clknet_leaf_66_wb_clk_i _02226_ _00461_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.ADR_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17431__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15549_ net1278 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09070_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[18\] net658 _05325_ _05328_
+ _05331_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_115_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ clknet_leaf_120_wb_clk_i _02779_ _01082_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_18199_ net1573 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
XFILLER_0_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17581__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__A1 _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[18\] vssd1 vssd1 vccd1 vccd1
+ net2329 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09087__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold724 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold746 team_01_WB.instance_to_wrap.cpu.RF0.registers\[7\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08422__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold757 team_01_WB.instance_to_wrap.cpu.RF0.registers\[26\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15817__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold768 _02039_ vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10026__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold779 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap487 _04344_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_1
X_09972_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[21\]\[5\] net619 _06217_ _06228_
+ _06230_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14721__A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14141__A2 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[21\] net617 _05170_ _05179_
+ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09815__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout297_A _08001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__C1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1402 team_01_WB.instance_to_wrap.cpu.FetchedInstr\[24\] vssd1 vssd1 vccd1 vccd1
+ net3018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net3029 sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ net1073 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[20\] net885
+ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and3_1
Xhold1424 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net3040 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1004_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1435 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net3051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1446 team_01_WB.instance_to_wrap.cpu.RF0.registers\[18\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net3062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08785_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[22\] net660 net650 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\]
+ _05048_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a221o_1
Xhold1457 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net3073
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 net3084
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09253__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1479 _03472_ vssd1 vssd1 vccd1 vccd1 net3095 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout464_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13101__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16529__CLK clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12387__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11663__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout631_A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1373_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ net1068 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[13\] net871
+ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09337_ net1000 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[14\] net896 vssd1
+ vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16679__CLK clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09268_ net1070 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[15\] net847
+ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[12\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[15\]
+ team_01_WB.instance_to_wrap.cpu.FetchedInstr\[14\] team_01_WB.instance_to_wrap.cpu.FetchedInstr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__or4b_1
XFILLER_0_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09199_ net1077 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[16\] net877
+ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13011__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12915__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11230_ net547 _07493_ _07491_ _07485_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09387__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09428__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _06319_ _06597_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12850__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10112_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[3\] _04765_ _06353_
+ _06354_ _06356_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14132__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _05993_ _05788_ net504 vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13340__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[31\]\[4\] net632 _06289_ _06293_
+ _06298_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17304__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14920_ net1208 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 team_01_WB.instance_to_wrap.cpu.RF0.registers\[0\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_01_WB.instance_to_wrap.cpu.f0.write_data\[5\] vssd1 vssd1 vccd1 vccd1
+ net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_01_WB.instance_to_wrap.cpu.f0.write_data\[22\] vssd1 vssd1 vccd1 vccd1
+ net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 team_01_WB.instance_to_wrap.cpu.f0.write_data\[17\] vssd1 vssd1 vccd1 vccd1
+ net1689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ net1353 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XANTENNA__09163__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 net1700
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_01_WB.instance_to_wrap.cpu.f0.write_data\[9\] vssd1 vssd1 vccd1 vccd1
+ net1711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _04476_ _07771_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17570_ clknet_leaf_143_wb_clk_i _03130_ _01433_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14782_ net1382 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XANTENNA__13643__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ net2853 net299 net468 vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
XANTENNA__11103__C1 _07363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10102__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16521_ clknet_leaf_73_wb_clk_i _02149_ _00384_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09311__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09460__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ team_01_WB.instance_to_wrap.cpu.f0.i\[24\] net1062 _07752_ _04025_ net485
+ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__o311a_1
XFILLER_0_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11654__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12297__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ _06697_ _06752_ _06807_ _04988_ net498 net514 vssd1 vssd1 vccd1 vccd1 _07209_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16452_ clknet_leaf_106_wb_clk_i net2076 _00315_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14199__A2 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13664_ net773 _07396_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10876_ net535 _07139_ _07138_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__o21ai_2
X_15403_ net1206 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12615_ net3017 net276 net397 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XANTENNA__11214__B _07477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16383_ clknet_leaf_82_wb_clk_i _00000_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13595_ net768 _07243_ net1067 vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18122_ net1496 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
X_15334_ net1274 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
X_12546_ net3010 net253 net405 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053_ net1615 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15265_ net1312 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
X_12477_ net1793 net285 net413 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
X_17004_ clknet_leaf_47_wb_clk_i _02564_ _00867_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12906__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 team_01_WB.instance_to_wrap.cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14216_ net1883 net585 net1171 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09378__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _07687_ net1626 _07685_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__mux2_1
XANTENNA__09338__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15196_ net1277 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11185__A2 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14147_ _04293_ _04298_ _04303_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__or4_1
XANTENNA__15637__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _05348_ _07224_ _05347_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__o21a_1
XANTENNA__18013__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[32\] _04238_ _04239_ team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[104\]
+ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13029_ net1717 net836 net355 _03672_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
X_17906_ clknet_leaf_78_wb_clk_i _03456_ _01726_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10145__B1 _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13882__A1 _04505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 team_01_WB.instance_to_wrap.cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1
+ net1060 sky130_fd_sc_hd__clkbuf_2
X_18202__1576 vssd1 vssd1 vccd1 vccd1 _18202__1576/HI net1576 sky130_fd_sc_hd__conb_1
XANTENNA__13882__B2 _07834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1071 net1105 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09550__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17837_ clknet_leaf_92_wb_clk_i _03388_ _01658_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.IM0.address_IM\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1082 net1088 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_1
Xfanout1093 net1096 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_1
XFILLER_0_94_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08570_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[30\] net660 net642 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a22o_1
X_17768_ clknet_leaf_97_wb_clk_i net1929 _01589_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.DM0.readdata\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09370__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16719_ clknet_leaf_54_wb_clk_i _02279_ _00582_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17699_ clknet_leaf_71_wb_clk_i _03259_ _01538_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.K0.code\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12000__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18130__1504 vssd1 vssd1 vccd1 vccd1 _18130__1504/HI net1504 sky130_fd_sc_hd__conb_1
XFILLER_0_92_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10852__A1_N net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09122_ net1011 team_01_WB.instance_to_wrap.cpu.RF0.registers\[15\]\[17\] net862
+ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ net1083 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[18\] net845
+ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold521 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08577__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _02030_ vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 team_01_WB.instance_to_wrap.cpu.c0.count\[4\] vssd1 vssd1 vccd1 vccd1 net2170
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12670__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17327__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 team_01_WB.instance_to_wrap.cpu.RF0.registers\[20\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10384__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_01_WB.instance_to_wrap.cpu.RF0.registers\[10\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold587 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11794__B _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 team_01_WB.instance_to_wrap.cpu.RF0.registers\[28\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[1\]\[5\] net852 vssd1
+ vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13322__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net1076 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[21\] net884
+ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__and3_1
XANTENNA__10136__B1 _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ net1023 team_01_WB.instance_to_wrap.cpu.RF0.registers\[6\]\[6\] net844 vssd1
+ vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__and3_1
Xhold1210 team_01_WB.instance_to_wrap.cpu.RF0.registers\[12\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_01_WB.instance_to_wrap.cpu.RF0.registers\[2\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 team_01_WB.instance_to_wrap.cpu.RF0.registers\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 team_01_WB.instance_to_wrap.cpu.LCD0.row_2\[105\] vssd1 vssd1 vccd1 vccd1
+ net2859 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net1010 team_01_WB.instance_to_wrap.cpu.RF0.registers\[11\]\[20\] net865
+ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1254 _02086_ vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1265 team_01_WB.instance_to_wrap.cpu.RF0.registers\[22\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15282__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1276 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 team_01_WB.instance_to_wrap.cpu.RF0.registers\[4\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ team_01_WB.instance_to_wrap.cpu.RF0.registers\[14\]\[22\] net738 net729 team_01_WB.instance_to_wrap.cpu.RF0.registers\[30\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09711__C net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08699_ net1118 team_01_WB.instance_to_wrap.cpu.RF0.registers\[24\]\[23\] net956
+ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13006__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11315__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ _06986_ _06993_ _06992_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__or3b_1
XFILLER_0_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10661_ _05481_ _05448_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12845__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ net2914 net196 net421 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__mux2_1
X_13380_ net2791 net326 net350 team_01_WB.instance_to_wrap.cpu.f0.i\[18\] vssd1 vssd1
+ vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10592_ _06849_ _06852_ _06855_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__or3_4
XFILLER_0_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ net3013 net211 net430 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12262_ net2140 net308 net437 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__mux2_1
X_15050_ net1220 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09158__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14001_ _04163_ _04179_ _04171_ _04167_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08568__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ _07107_ _07474_ _07476_ _07469_ _06315_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12580__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ net2143 net299 net446 vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
XANTENNA__12903__A3 _03605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08997__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11144_ _07248_ _07407_ net523 vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__mux2_1
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15952_ net1330 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__inv_2
X_11075_ _07087_ _07114_ net523 vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10026_ net1019 team_01_WB.instance_to_wrap.cpu.RF0.registers\[5\]\[4\] net859 vssd1
+ vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and3_1
X_14903_ net1257 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
X_15883_ net1352 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__inv_2
XANTENNA__11924__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ clknet_leaf_33_wb_clk_i _03182_ _01485_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13705__A team_01_WB.instance_to_wrap.cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14834_ net1343 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13616__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09190__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17553_ clknet_leaf_22_wb_clk_i _03113_ _01416_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14765_ net1189 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XANTENNA__13092__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11977_ net3252 net198 net467 vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ clknet_leaf_106_wb_clk_i _02132_ _00367_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[116\]
+ sky130_fd_sc_hd__dfstp_1
X_13716_ team_01_WB.instance_to_wrap.cpu.f0.i\[27\] _04021_ vssd1 vssd1 vccd1 vccd1
+ _04036_ sky130_fd_sc_hd__nand2_1
X_17484_ clknet_leaf_44_wb_clk_i _03044_ _01347_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.RF0.registers\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10928_ _05203_ net339 _07190_ _07191_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14696_ net1405 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16435_ clknet_leaf_101_wb_clk_i net1733 _00298_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.cpu.LCD0.row_1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10850__A1 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12755__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ net769 _07510_ net1067 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ _06830_ _07122_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16366_ clknet_leaf_66_wb_clk_i net1968 _00234_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08534__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13578_ _03902_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18105_ net1479 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
X_15317_ net1173 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XANTENNA__16224__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ net2225 net290 net409 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16297_ clknet_leaf_111_wb_clk_i _01931_ _00165_ vssd1 vssd1 vccd1 vccd1 team_01_WB.instance_to_wrap.a1.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18036_ net1602 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_15248_ net1262 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
XANTENNA__09068__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08559__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12490__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ net1205 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16374__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net310 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_0_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08700__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ net1005 team_01_WB.instance_to_wrap.cpu.RF0.registers\[9\]\[10\] net891 vssd1
+ vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and3_1
XANTENNA__10304__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

