`default_nettype none
module t06_lcd1602 (
	clk,
	rst,
	row_1,
	row_2,
	lcd_en,
	lcd_rw,
	lcd_rs,
	lcd_data
);
	parameter clk_div = 24000;
	input clk;
	input rst;
	input [127:0] row_1;
	input [127:0] row_2;
	output wire lcd_en;
	output wire lcd_rw;
	output reg lcd_rs;
	output reg [7:0] lcd_data;
	wire lcd_ctrl;
	reg [7:0] currentState;
	reg [7:0] nextState;
	reg [17:0] cnt_20ms;
	reg [14:0] cnt_500hz;
	wire delay_done;
	localparam TIME_500HZ = clk_div;
	localparam TIME_20MS = TIME_500HZ * 10;
	localparam IDLE_LCD = 8'h00;
	localparam SET_FUNCTION = 8'h01;
	localparam DISP_OFF = 8'h03;
	localparam DISP_CLEAR = 8'h02;
	localparam ENTRY_MODE = 8'h06;
	localparam DISP_ON = 8'h07;
	localparam ROW1_ADDR = 8'h05;
	localparam ROW1_0 = 8'h04;
	localparam ROW1_1 = 8'h0c;
	localparam ROW1_2 = 8'h0d;
	localparam ROW1_3 = 8'h0f;
	localparam ROW1_4 = 8'h0e;
	localparam ROW1_5 = 8'h0a;
	localparam ROW1_6 = 8'h0b;
	localparam ROW1_7 = 8'h09;
	localparam ROW1_8 = 8'h08;
	localparam ROW1_9 = 8'h18;
	localparam ROW1_A = 8'h19;
	localparam ROW1_B = 8'h1b;
	localparam ROW1_C = 8'h1a;
	localparam ROW1_D = 8'h1e;
	localparam ROW1_E = 8'h1f;
	localparam ROW1_F = 8'h1d;
	localparam ROW2_ADDR = 8'h1c;
	localparam ROW2_0 = 8'h14;
	localparam ROW2_1 = 8'h15;
	localparam ROW2_2 = 8'h17;
	localparam ROW2_3 = 8'h16;
	localparam ROW2_4 = 8'h12;
	localparam ROW2_5 = 8'h13;
	localparam ROW2_6 = 8'h11;
	localparam ROW2_7 = 8'h10;
	localparam ROW2_8 = 8'h30;
	localparam ROW2_9 = 8'h31;
	localparam ROW2_A = 8'h33;
	localparam ROW2_B = 8'h32;
	localparam ROW2_C = 8'h36;
	localparam ROW2_D = 8'h37;
	localparam ROW2_E = 8'h35;
	localparam ROW2_F = 8'h34;
	assign delay_done = (cnt_20ms == (TIME_20MS - 1) ? 1'b1 : 1'b0);
	always @(posedge clk)
		if (!rst)
			cnt_20ms <= 0;
		else if (cnt_20ms == (TIME_20MS - 1))
			cnt_20ms <= cnt_20ms;
		else
			cnt_20ms <= cnt_20ms + 1;
	always @(posedge clk)
		if (!rst)
			cnt_500hz <= 0;
		else if (delay_done) begin
			if (cnt_500hz == (TIME_500HZ - 1))
				cnt_500hz <= 0;
			else
				cnt_500hz <= cnt_500hz + 1;
		end
		else
			cnt_500hz <= 0;
	assign lcd_en = (cnt_500hz > ((TIME_500HZ - 1) / 2) ? 1'b0 : 1'b1);
	assign lcd_ctrl = (cnt_500hz == (TIME_500HZ - 1) ? 1'b1 : 1'b0);
	always @(posedge clk)
		if (!rst)
			currentState <= IDLE_LCD;
		else if (lcd_ctrl)
			currentState <= nextState;
		else
			currentState <= currentState;
	always @(*)
		case (currentState)
			IDLE_LCD: nextState = SET_FUNCTION;
			SET_FUNCTION: nextState = DISP_OFF;
			DISP_OFF: nextState = DISP_CLEAR;
			DISP_CLEAR: nextState = ENTRY_MODE;
			ENTRY_MODE: nextState = DISP_ON;
			DISP_ON: nextState = ROW1_ADDR;
			ROW1_ADDR: nextState = ROW1_0;
			ROW1_0: nextState = ROW1_1;
			ROW1_1: nextState = ROW1_2;
			ROW1_2: nextState = ROW1_3;
			ROW1_3: nextState = ROW1_4;
			ROW1_4: nextState = ROW1_5;
			ROW1_5: nextState = ROW1_6;
			ROW1_6: nextState = ROW1_7;
			ROW1_7: nextState = ROW1_8;
			ROW1_8: nextState = ROW1_9;
			ROW1_9: nextState = ROW1_A;
			ROW1_A: nextState = ROW1_B;
			ROW1_B: nextState = ROW1_C;
			ROW1_C: nextState = ROW1_D;
			ROW1_D: nextState = ROW1_E;
			ROW1_E: nextState = ROW1_F;
			ROW1_F: nextState = ROW2_ADDR;
			ROW2_ADDR: nextState = ROW2_0;
			ROW2_0: nextState = ROW2_1;
			ROW2_1: nextState = ROW2_2;
			ROW2_2: nextState = ROW2_3;
			ROW2_3: nextState = ROW2_4;
			ROW2_4: nextState = ROW2_5;
			ROW2_5: nextState = ROW2_6;
			ROW2_6: nextState = ROW2_7;
			ROW2_7: nextState = ROW2_8;
			ROW2_8: nextState = ROW2_9;
			ROW2_9: nextState = ROW2_A;
			ROW2_A: nextState = ROW2_B;
			ROW2_B: nextState = ROW2_C;
			ROW2_C: nextState = ROW2_D;
			ROW2_D: nextState = ROW2_E;
			ROW2_E: nextState = ROW2_F;
			ROW2_F: nextState = ROW1_ADDR;
			default: nextState = IDLE_LCD;
		endcase
	assign lcd_rw = 1'b0;
	always @(posedge clk)
		if (!rst)
			lcd_rs <= 1'b0;
		else if (lcd_ctrl) begin
			if (((((((nextState == SET_FUNCTION) || (nextState == DISP_OFF)) || (nextState == DISP_CLEAR)) || (nextState == ENTRY_MODE)) || (nextState == DISP_ON)) || (nextState == ROW1_ADDR)) || (nextState == ROW2_ADDR))
				lcd_rs <= 1'b0;
			else
				lcd_rs <= 1'b1;
		end
		else
			lcd_rs <= lcd_rs;
	always @(posedge clk)
		if (!rst)
			lcd_data <= 8'h00;
		else if (lcd_ctrl)
			case (nextState)
				IDLE_LCD: lcd_data <= 8'hxx;
				SET_FUNCTION: lcd_data <= 8'h38;
				DISP_OFF: lcd_data <= 8'h08;
				DISP_CLEAR: lcd_data <= 8'h01;
				ENTRY_MODE: lcd_data <= 8'h06;
				DISP_ON: lcd_data <= 8'h0c;
				ROW1_ADDR: lcd_data <= 8'h80;
				ROW1_0: lcd_data <= row_1[127:120];
				ROW1_1: lcd_data <= row_1[119:112];
				ROW1_2: lcd_data <= row_1[111:104];
				ROW1_3: lcd_data <= row_1[103:96];
				ROW1_4: lcd_data <= row_1[95:88];
				ROW1_5: lcd_data <= row_1[87:80];
				ROW1_6: lcd_data <= row_1[79:72];
				ROW1_7: lcd_data <= row_1[71:64];
				ROW1_8: lcd_data <= row_1[63:56];
				ROW1_9: lcd_data <= row_1[55:48];
				ROW1_A: lcd_data <= row_1[47:40];
				ROW1_B: lcd_data <= row_1[39:32];
				ROW1_C: lcd_data <= row_1[31:24];
				ROW1_D: lcd_data <= row_1[23:16];
				ROW1_E: lcd_data <= row_1[15:8];
				ROW1_F: lcd_data <= row_1[7:0];
				ROW2_ADDR: lcd_data <= 8'hc0;
				ROW2_0: lcd_data <= row_2[127:120];
				ROW2_1: lcd_data <= row_2[119:112];
				ROW2_2: lcd_data <= row_2[111:104];
				ROW2_3: lcd_data <= row_2[103:96];
				ROW2_4: lcd_data <= row_2[95:88];
				ROW2_5: lcd_data <= row_2[87:80];
				ROW2_6: lcd_data <= row_2[79:72];
				ROW2_7: lcd_data <= row_2[71:64];
				ROW2_8: lcd_data <= row_2[63:56];
				ROW2_9: lcd_data <= row_2[55:48];
				ROW2_A: lcd_data <= row_2[47:40];
				ROW2_B: lcd_data <= row_2[39:32];
				ROW2_C: lcd_data <= row_2[31:24];
				ROW2_D: lcd_data <= row_2[23:16];
				ROW2_E: lcd_data <= row_2[15:8];
				ROW2_F: lcd_data <= row_2[7:0];
				default: lcd_data <= 8'hxx;
			endcase
		else
			lcd_data <= lcd_data;
endmodule
