* NGSPICE file created from team_02.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_02 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8]
+ gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14]
+ gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20]
+ gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27]
+ gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[3] gpio_oeb[4]
+ gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10]
+ gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17]
+ gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23]
+ gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2]
+ gpio_out[30] gpio_out[31] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XPHY_EDGE_ROW_176_Left_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06883_ top.DUT.register\[2\]\[22\] net717 net699 top.DUT.register\[23\]\[22\] _02009_
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a221o_1
X_09671_ _03353_ net340 net336 _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_124_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08622_ net890 top.pc\[15\] net539 _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a22o_1
X_08553_ net886 top.pc\[12\] net537 _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07504_ net809 net498 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08484_ _02235_ net469 _03599_ net520 _03600_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o221a_1
XANTENNA__07837__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07435_ _02555_ _02561_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__nor2_4
XANTENNA__09039__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_185_Left_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1071_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07366_ net499 _02492_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__or2_2
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06317_ _01451_ _01332_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__and2_1
X_09105_ _01587_ _04162_ _04163_ _01614_ _04049_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a32o_1
XANTENNA__10185__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ top.a1.instruction\[21\] net524 _01621_ top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 _02424_ sky130_fd_sc_hd__a22o_1
XANTENNA__06207__C_N net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09036_ net321 _03374_ _03448_ _03744_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a211o_1
XANTENNA__09974__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06248_ net1469 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[24\] sky130_fd_sc_hd__and2_1
XANTENNA__07470__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 top.DUT.register\[27\]\[25\] vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ net913 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
XANTENNA__10913__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 top.DUT.register\[4\]\[25\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 top.DUT.register\[29\]\[21\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold373 top.DUT.register\[28\]\[0\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 top.DUT.register\[11\]\[12\] vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 top.ramaddr\[14\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 _05022_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_2
Xfanout842 _05023_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_2
X_09938_ net223 net2164 net433 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__mux2_1
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_2
Xfanout864 _01430_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_4
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_181_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout886 net889 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _04543_ net527 net333 top.a1.dataIn\[26\] net335 vssd1 vssd1 vccd1 vccd1
+ _04866_ sky130_fd_sc_hd__a221o_1
Xfanout897 net899 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__clkbuf_4
Xhold1040 top.DUT.register\[10\]\[11\] vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 top.DUT.register\[7\]\[11\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1062 top.pad.button_control.r_counter\[7\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ _05733_ _05750_ _05768_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1073 top.DUT.register\[15\]\[17\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ clknet_leaf_0_clk _00444_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1084 top.DUT.register\[8\]\[19\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 top.DUT.register\[3\]\[27\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11831_ _05653_ _05654_ _05677_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__and3_1
XANTENNA__09278__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07289__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ _05598_ _05631_ _05604_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12603__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13501_ clknet_leaf_103_clk _01065_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ net244 net1676 net383 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
X_11693_ _05552_ _05556_ _05557_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13432_ clknet_leaf_109_clk _00996_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ net1391 net265 net451 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09045__A4 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575_ net158 net2110 net359 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
X_13363_ clknet_leaf_5_clk _00927_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10095__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09884__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ top.lcd.cnt_500hz\[12\] _06114_ _06116_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__o21a_1
X_13294_ clknet_leaf_117_clk _00858_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12245_ top.lcd.cnt_20ms\[3\] _06063_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__xor2_1
XANTENNA__10823__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08005__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07213__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ _06019_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07764__A1 _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11127_ net55 net857 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and2_1
XFILLER_0_208_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ net104 net860 net829 net1190 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08713__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ net208 net2203 net426 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07220_ top.DUT.register\[21\]\[15\] net573 net571 top.DUT.register\[8\]\[15\] _02346_
+ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07151_ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07082_ top.a1.instruction\[7\] _01477_ _01620_ top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 _02209_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_89_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10733__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09095__A _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07755__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06558__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08952__B1 _02757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout127 _05878_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_2
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout149 _04691_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_1
X_07984_ top.DUT.register\[12\]\[31\] net582 net745 top.DUT.register\[31\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__a22o_1
X_09723_ net894 net534 _04318_ net823 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a31o_1
X_06935_ top.DUT.register\[30\]\[21\] net618 _02061_ vssd1 vssd1 vccd1 vccd1 _02062_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout377_A _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__B1 _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ top.a1.instruction\[11\] _04675_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__nand2_1
X_06866_ _01973_ _01991_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08605_ _02361_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _04615_ _04616_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a21oi_1
X_06797_ top.DUT.register\[22\]\[24\] net754 net727 top.DUT.register\[10\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout544_A _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06730__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09969__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ _03456_ _03650_ net310 vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_193_Left_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07630__X _02757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08467_ net321 _03545_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10908__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09680__A1 top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07418_ top.DUT.register\[14\]\[6\] net722 net707 top.DUT.register\[15\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07691__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08398_ net476 _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__or2_1
Xwire517 _01885_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07349_ top.DUT.register\[21\]\[8\] net572 net639 top.DUT.register\[11\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a22o_1
XANTENNA__11312__B top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07443__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10360_ net1450 net176 net393 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06797__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ _03456_ _03537_ net273 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a21o_1
X_10291_ net1570 net184 net404 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
XANTENNA__10643__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _05886_ _05888_ _05894_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nor4_1
Xhold170 top.ramaddr\[6\] vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 top.a1.row1\[115\] vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06549__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 top.a1.row1\[109\] vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout650 _01642_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_4
Xfanout672 net673 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_8
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ clknet_leaf_40_clk _00496_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12863_ clknet_leaf_115_clk _00427_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ _05682_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12794_ clknet_leaf_16_clk _00358_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _05589_ _05600_ _05593_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09671__A1 _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10818__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _05544_ _05545_ _05542_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13415_ clknet_leaf_25_clk _00979_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10627_ net230 net2148 net390 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__mux2_1
XANTENNA__09423__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13346_ clknet_leaf_42_clk _00910_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10558_ net221 net2204 net359 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10553__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ clknet_leaf_107_clk _00841_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10489_ net235 net2241 net365 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__mux2_1
X_12228_ _05984_ net589 _06062_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _06024_ _06025_ _06027_ _06022_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_208_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06960__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12596__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ top.DUT.register\[13\]\[26\] net649 net565 top.DUT.register\[4\]\[26\] _01846_
+ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a221o_1
XANTENNA__09362__B _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12525__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire512_A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06651_ _01776_ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__nor2_2
XANTENNA__09074__D_N _02685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13869__1156 vssd1 vssd1 vccd1 vccd1 net1156 _13869__1156/LO sky130_fd_sc_hd__conb_1
X_09370_ _04413_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or2_1
X_06582_ top.DUT.register\[17\]\[29\] net724 net679 top.DUT.register\[13\]\[29\] _01708_
+ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08321_ net311 _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10728__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ _02883_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07673__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ top.DUT.register\[9\]\[15\] net708 net667 top.DUT.register\[5\]\[15\] _02321_
+ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08183_ _03307_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07134_ top.DUT.register\[28\]\[12\] net653 net605 top.DUT.register\[18\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a22o_1
XANTENNA__07425__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08968__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07065_ net794 _02190_ _02191_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__or3b_1
XANTENNA__10463__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1034_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07728__A1 _02854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _01994_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout759_A _01510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07344__Y _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ net836 _04256_ _04720_ top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 _04721_
+ sky130_fd_sc_hd__a2bb2o_1
X_06918_ top.DUT.register\[5\]\[21\] net670 _02042_ _02044_ vssd1 vssd1 vccd1 vccd1
+ _02045_ sky130_fd_sc_hd__a211o_1
X_07898_ top.DUT.register\[21\]\[17\] net572 net560 top.DUT.register\[23\]\[17\] _03024_
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a221o_1
XANTENNA__09840__X _04840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09637_ _04645_ _04646_ _01472_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__o21ai_1
X_06849_ top.DUT.register\[12\]\[23\] net580 net739 top.DUT.register\[8\]\[23\] _01975_
+ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout926_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ top.pc\[29\] top.pc\[30\] _04566_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08519_ _02164_ net483 net469 _02165_ _03627_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__o221a_1
XFILLER_0_194_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10638__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ top.pc\[26\] _04518_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07664__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ _05341_ _05363_ _05369_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__or3b_1
XFILLER_0_25_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ _05289_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13200_ clknet_leaf_0_clk _00764_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10412_ net144 net1720 net328 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11392_ _05236_ _05256_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ clknet_leaf_30_clk _00695_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10343_ net1642 net243 net394 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XANTENNA__09708__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net1560 net246 net401 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__mux2_1
X_13062_ clknet_leaf_19_clk _00626_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12013_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__inv_2
XANTENNA__08392__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__A2 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__B2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09463__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06942__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout480 _03255_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08079__A _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ clknet_leaf_1_clk _00479_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11217__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09892__B2 top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ clknet_leaf_116_clk _00410_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ clknet_leaf_2_clk _00341_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10548__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ top.a1.dataIn\[10\] _05526_ _05527_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_211_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07407__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold906 top.DUT.register\[20\]\[26\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07958__A1 _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold917 top.DUT.register\[2\]\[27\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ clknet_leaf_110_clk _00893_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10283__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold928 top.DUT.register\[15\]\[29\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 top.DUT.register\[31\]\[11\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_08870_ net478 _03964_ _03968_ net481 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07186__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07821_ net806 _02947_ _01624_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06933__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07752_ _02877_ _02878_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__and2b_1
XANTENNA__07605__B _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06703_ top.DUT.register\[25\]\[26\] net773 net750 top.DUT.register\[20\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11127__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ net805 _02788_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09883__A1 _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A2 top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _04459_ _04463_ _01619_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__a21o_1
X_06634_ top.DUT.register\[9\]\[28\] net629 net601 top.DUT.register\[10\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a22o_1
XANTENNA__07894__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10966__B net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ net132 _04392_ _04399_ net819 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__o22a_1
XANTENNA__09635__A1 top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10458__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06565_ _01560_ _01690_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout242_A _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08304_ _03177_ _03414_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07646__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06496_ top.a1.instruction\[31\] _01622_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__nand2_2
X_09284_ top.pc\[13\] _04318_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__xor2_1
XANTENNA__07110__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08235_ net276 _03229_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08166_ net286 _03291_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07117_ top.DUT.register\[4\]\[12\] net770 _01520_ top.DUT.register\[17\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
X_08097_ net495 net295 vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10193__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06204__A_N top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09267__B _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09982__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload90 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__07068__A _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ _02167_ _02171_ _02172_ _02174_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__or4_2
XANTENNA__10921__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12447__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _03942_ _03960_ _04060_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__and3_1
XANTENNA__06924__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10961_ top.a1.halfData\[5\] _01413_ _01415_ _01381_ _01410_ vssd1 vssd1 vccd1 vccd1
+ _04987_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_3_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_206_Right_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ clknet_leaf_53_clk _00264_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09730__B _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ clknet_leaf_94_clk _00012_ net993 vssd1 vssd1 vccd1 vccd1 top.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10892_ net2301 net184 net348 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ clknet_leaf_106_clk _00195_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12149__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07637__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12562_ clknet_leaf_51_clk _00126_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07101__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ _05349_ _05371_ _05353_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ clknet_leaf_82_clk _00060_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramstore\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11444_ _05277_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11375_ _05214_ _05239_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09714__A1_N net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13114_ clknet_leaf_18_clk _00678_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ net2338 net175 net397 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
X_13868__1155 vssd1 vssd1 vccd1 vccd1 net1155 _13868__1155/LO sky130_fd_sc_hd__conb_1
Xclkbuf_4_2__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_13045_ clknet_leaf_8_clk _00609_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08970__A1_N _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ net1483 net176 net454 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__mux2_1
XANTENNA__10831__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07168__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ net187 net1933 net411 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
XANTENNA__06915__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08668__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07876__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ net1129 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__08537__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07340__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ clknet_leaf_112_clk _00393_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10278__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06350_ net34 top.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__nand2_1
XANTENNA__07628__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06281_ net1497 net878 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[25\] sky130_fd_sc_hd__and2_1
XFILLER_0_44_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ net808 _03146_ net463 vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__o21a_1
XANTENNA__09368__A top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 top.DUT.register\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 top.DUT.register\[2\]\[6\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold725 top.DUT.register\[26\]\[25\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 top.DUT.register\[27\]\[28\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 top.DUT.register\[8\]\[18\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 top.DUT.register\[28\]\[20\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ net1673 net231 net430 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
Xhold769 top.DUT.register\[9\]\[24\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ _03107_ _03152_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10741__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07159__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__RESET_B net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ net482 _03949_ _03950_ net520 _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout192_A _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07804_ top.DUT.register\[16\]\[19\] net637 net547 top.DUT.register\[5\]\[19\] _02930_
+ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a221o_1
X_08784_ net305 _03823_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08108__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A_N _02298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07735_ top.DUT.register\[22\]\[1\] net754 net741 top.DUT.register\[8\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a22o_1
XANTENNA__10977__A top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07666_ top.DUT.register\[17\]\[0\] net643 net635 top.DUT.register\[16\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07331__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13327__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _04446_ _04447_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__nor2_1
X_06617_ top.DUT.register\[22\]\[28\] net753 net733 top.DUT.register\[19\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a22o_1
XANTENNA__10188__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ _02715_ _02717_ _02721_ _02723_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout624_A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07619__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ net819 _04383_ _04377_ _04186_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_173_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06548_ top.DUT.register\[17\]\[30\] net644 net620 top.DUT.register\[26\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ net507 _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10916__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06479_ net902 _01388_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11601__A top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ net476 _03332_ net469 _02880_ _03337_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__o221a_1
XFILLER_0_160_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08182__A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ top.pc\[8\] _04241_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08149_ net297 _03012_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07398__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ top.a1.data\[2\] net797 _05000_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ net1323 net200 net460 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
XANTENNA__10651__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11091_ net67 net858 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ net220 net1705 net424 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__mux2_1
Xhold30 top.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 top.a1.data\[10\] vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 net116 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 _01189_ vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold74 _01198_ vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 top.ramaddr\[30\] vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_65_clk _01344_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07570__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold96 top.ramstore\[16\] vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _05836_ _05846_ _05837_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o21a_1
Xclkbuf_4_10__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13732_ clknet_leaf_73_clk _01275_ net1091 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07858__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ _04628_ net847 vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_67_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13663_ clknet_leaf_88_clk _01222_ net1005 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
X_10875_ net1819 net246 net345 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12614_ clknet_leaf_23_clk _00178_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ clknet_leaf_97_clk _01153_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12545_ clknet_leaf_80_clk _00109_ net1002 vssd1 vssd1 vccd1 vccd1 top.pc\[28\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10826__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12476_ clknet_leaf_95_clk top.ru.next_FetchedInstr\[28\] net991 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[28\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11230__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _05295_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__or2_1
XANTENNA_5 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__B1 _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08586__A1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _05199_ _05227_ _05197_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06597__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net2067 net245 net399 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XANTENNA__10561__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ top.a1.row1\[108\] _05161_ _05164_ _05156_ _05160_ vssd1 vssd1 vccd1 vccd1
+ _05165_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_169_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08338__B2 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ clknet_leaf_40_clk _00592_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_206_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1050 net1051 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1063 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
Xfanout1072 net1076 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_2
XFILLER_0_177_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1083 net1084 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
Xfanout1094 net1097 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09299__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ top.DUT.register\[1\]\[4\] net657 net626 top.DUT.register\[25\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XANTENNA__07849__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07313__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07171__A _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12785__Q top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07451_ top.DUT.register\[23\]\[6\] net562 net638 top.DUT.register\[16\]\[6\] _02577_
+ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06402_ _01496_ _01499_ net791 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07382_ top.DUT.register\[25\]\[7\] net772 net736 top.DUT.register\[24\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09121_ net895 top.pc\[3\] vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__nand2_1
X_06333_ _01449_ _01470_ _01471_ _01334_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _03433_ _04069_ _04112_ _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__and4_1
X_06264_ net1829 net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[8\] sky130_fd_sc_hd__and2_1
XFILLER_0_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09098__A _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08003_ top.DUT.register\[13\]\[31\] net649 net597 top.DUT.register\[27\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a22o_1
X_06195_ top.a1.halfData\[0\] _01411_ _01415_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__and3_1
Xhold500 top.DUT.register\[27\]\[27\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 top.DUT.register\[16\]\[1\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 top.DUT.register\[19\]\[8\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 top.DUT.register\[16\]\[13\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold544 top.DUT.register\[23\]\[11\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 top.DUT.register\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 top.DUT.register\[21\]\[26\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 top.lcd.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 top.DUT.register\[10\]\[8\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10471__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09954_ net166 net1696 net435 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__mux2_1
Xhold599 top.DUT.register\[19\]\[18\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ net305 _03929_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10136__A1 top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _03973_ net343 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout574_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08836_ _01862_ net484 _03936_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07552__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__X _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08767_ net272 _03725_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__nand2_1
XANTENNA__09829__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06760__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07718_ top.DUT.register\[28\]\[1\] net653 net625 top.DUT.register\[25\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__a22o_1
X_08698_ net271 _03624_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07304__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07081__A top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07649_ top.DUT.register\[25\]\[2\] net771 net751 top.DUT.register\[22\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867__1154 vssd1 vssd1 vccd1 vccd1 net1154 _13867__1154/LO sky130_fd_sc_hd__conb_1
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ net2106 net217 net450 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12867__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ net135 _04360_ _04367_ net819 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_62_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10646__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_114_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10591_ net207 net1535 net388 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XANTENNA__10072__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[2\]
+ top.pad.button_control.r_counter\[1\] vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08017__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net1249 _06082_ _06084_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__a21oi_1
X_11212_ net882 net884 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_186_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12192_ net1343 net846 net814 _06059_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06579__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
X_11143_ net64 net859 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and2_1
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07791__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__clkbuf_4
X_11074_ net90 net856 net825 net1258 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ net158 net1966 net427 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
XANTENNA__07543__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08358__Y _03480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _05825_ _05845_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_88_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13715_ clknet_leaf_71_clk _01263_ net1096 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ net172 net1644 net444 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13646_ clknet_leaf_84_clk _01205_ net1015 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
X_10858_ net1522 net189 net351 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08815__A _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08256__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13577_ clknet_leaf_96_clk _01136_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_105_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10556__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10789_ net1685 net214 net448 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12528_ clknet_leaf_82_clk _00092_ net1013 vssd1 vssd1 vccd1 vccd1 top.pc\[11\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__11260__C1 _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08008__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ clknet_leaf_98_clk top.ru.next_FetchedInstr\[11\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[11\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10291__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 _02759_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13172__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _02056_ _02076_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__and2_1
X_09670_ top.a1.dataIn\[1\] net794 _04689_ top.pc\[1\] net343 vssd1 vssd1 vccd1 vccd1
+ _04692_ sky130_fd_sc_hd__a221o_1
X_06882_ top.DUT.register\[19\]\[22\] net733 net725 top.DUT.register\[17\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08621_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06742__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08552_ net473 _03645_ _03666_ net477 _03661_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07105__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07503_ _02614_ _02617_ _02628_ _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__nor4_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11135__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08483_ _02234_ _03177_ net483 _02233_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout155_A _04900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07434_ _02544_ _02545_ _02558_ _02560_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__or4_2
XFILLER_0_91_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10466__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07365_ _02471_ _02491_ net805 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _01589_ _04153_ _04165_ net833 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__and4b_1
X_06316_ _01450_ _01454_ _01455_ _01458_ _01449_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07296_ _02413_ _02417_ _02422_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__nor3_2
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08262__A3 _03386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09035_ net321 _03297_ _03744_ _04068_ _04076_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06247_ net1424 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[23\] sky130_fd_sc_hd__and2_1
XFILLER_0_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold330 top.DUT.register\[5\]\[1\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08460__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06178_ net36 net35 net38 net37 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__nor4_1
XANTENNA__06532__X _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 top.DUT.register\[12\]\[0\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 top.DUT.register\[28\]\[23\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 top.DUT.register\[11\]\[27\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 top.DUT.register\[14\]\[28\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold385 top.DUT.register\[14\]\[15\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 top.DUT.register\[30\]\[23\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout810 _01495_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
Xfanout832 _05022_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__dlymetal6s2s_1
X_09937_ net231 net1785 net434 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__mux2_1
Xfanout843 _04966_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06981__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_2
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout876 net878 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_2
X_09868_ net833 _04534_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nor2_1
Xfanout887 net889 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
Xhold1030 top.DUT.register\[21\]\[23\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08722__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1041 top.DUT.register\[12\]\[17\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1052 top.DUT.register\[20\]\[6\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08722__B2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ _01908_ _01950_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nor2_1
Xhold1063 top.DUT.register\[23\]\[28\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 top.DUT.register\[16\]\[20\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ net204 net1698 net439 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__mux2_1
Xhold1085 top.DUT.register\[5\]\[8\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11326__A top.a1.dataIn\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ _05672_ _05676_ _05652_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__a21o_1
Xhold1096 top.DUT.register\[4\]\[7\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11761_ _05589_ _05600_ _05595_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13500_ clknet_leaf_77_clk _01064_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10712_ net248 net1947 net382 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
X_11692_ _05556_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_3__f_clk_X clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13431_ clknet_leaf_77_clk _00995_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ net2003 net148 net450 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ clknet_leaf_51_clk _00926_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06155__A top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10574_ net162 net2285 net357 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ top.lcd.cnt_500hz\[12\] _06114_ net588 vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13293_ clknet_leaf_33_clk _00857_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08641__Y _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09738__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ _06071_ _06074_ net1108 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__o21a_1
XANTENNA__09466__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06442__X _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08410__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _06041_ _06044_ _06039_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07764__A2 _02586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11126_ net916 net1279 net853 _05049_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a31o_1
X_11057_ net103 net856 net825 net1183 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13431__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ net222 top.DUT.register\[4\]\[11\] net427 vssd1 vssd1 vccd1 vccd1 _00229_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output49_A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06724__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11236__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11959_ _05822_ _05823_ _05801_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08477__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13629_ clknet_leaf_61_clk net1285 net1100 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10286__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ _02275_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09441__A2 top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07081_ top.a1.instruction\[30\] _01621_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09095__B net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07755__A2 _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13866__1153 vssd1 vssd1 vccd1 vccd1 net1153 _13866__1153/LO sky130_fd_sc_hd__conb_1
XANTENNA__08952__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14__f_clk_X clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout139 _04181_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_07983_ top.DUT.register\[27\]\[31\] net777 net687 top.DUT.register\[1\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__a22o_1
XANTENNA__06963__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ net894 _01613_ _04318_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a21oi_1
X_06934_ top.DUT.register\[9\]\[21\] net629 net610 top.DUT.register\[12\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XANTENNA__13172__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09653_ top.a1.instruction\[11\] _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__and2_4
X_06865_ _01973_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__nor2_1
XANTENNA__06715__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _02401_ _03709_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__nand2_1
X_09584_ _04615_ _04616_ _01618_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o21ai_1
X_06796_ top.DUT.register\[28\]\[24\] net586 _01921_ _01922_ vssd1 vssd1 vccd1 vccd1
+ _01923_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ _03649_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout537_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ net317 _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__nor2_2
XFILLER_0_175_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ top.DUT.register\[22\]\[6\] net754 net745 top.DUT.register\[31\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10196__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_A _01533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _03516_ _03517_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire518 _01773_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_2
XANTENNA__09985__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ top.DUT.register\[17\]\[8\] net643 net607 top.DUT.register\[12\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10924__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07279_ top.DUT.register\[29\]\[9\] net701 net671 top.DUT.register\[16\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ _03683_ _03704_ net322 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07994__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10290_ net1480 net187 net404 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 top.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 top.ramaddr\[29\] vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 top.ramaddr\[25\] vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold193 top.a1.row1\[114\] vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06954__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _01648_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 _01641_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_8
Xfanout662 _01638_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout673 _01553_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_6
Xfanout684 _01544_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout695 _01540_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_8
X_12931_ clknet_leaf_33_clk _00495_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07534__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ clknet_leaf_13_clk _00426_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11813_ top.a1.dataIn\[7\] _05672_ _05676_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__and3_1
XANTENNA__12895__RESET_B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11058__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ clknet_leaf_36_clk _00357_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_194_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _05610_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__nor2_1
XANTENNA__07131__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09671__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11675_ _05512_ _05513_ _05541_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__and3_1
XANTENNA__09408__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13414_ clknet_leaf_24_clk _00978_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net179 top.DUT.register\[22\]\[15\] net389 vssd1 vssd1 vccd1 vccd1 _00809_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09748__X _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13345_ clknet_leaf_28_clk _00909_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12585__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ net225 net1600 net357 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__mux2_1
XANTENNA__10834__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09908__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ clknet_leaf_54_clk _00840_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10488_ net240 net1547 net366 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__mux2_1
X_12227_ net1238 net589 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nor2_1
XANTENNA__07198__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07737__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ _06022_ _06027_ _06026_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06945__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11109_ net45 net857 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_16_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12089_ _05949_ _05952_ _05953_ _05957_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__or4b_2
XFILLER_0_182_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06650_ _01755_ _01774_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__and2_1
XFILLER_0_189_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire505_A _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11049__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06581_ top.DUT.register\[25\]\[29\] net774 net695 top.DUT.register\[21\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ _03197_ _03211_ net302 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_50_clk_X clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07122__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08251_ _02783_ _02882_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08870__B1 _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07202_ top.DUT.register\[8\]\[15\] net740 net696 top.DUT.register\[23\]\[15\] _02326_
+ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a221o_1
XANTENNA_wire495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _02184_ net292 vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_41_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07133_ top.DUT.register\[29\]\[12\] net663 net554 top.DUT.register\[7\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08622__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10744__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07064_ net901 _01478_ _01577_ _01571_ _01481_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10980__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08492__A2_N _03606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1027_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06936__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__B _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _02015_ _02034_ _03092_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a21o_1
X_09705_ _04719_ _04716_ net534 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__mux2_4
X_06917_ top.DUT.register\[12\]\[21\] net583 net722 top.DUT.register\[14\]\[21\] _02043_
+ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ top.DUT.register\[17\]\[17\] net643 net595 top.DUT.register\[27\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_A _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09636_ _04644_ _04645_ _04646_ _04643_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o22ai_1
X_06848_ top.DUT.register\[26\]\[23\] net759 net704 top.DUT.register\[15\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a22o_1
XANTENNA__08737__X _03843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07361__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07900__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ _04595_ _04601_ top.pc\[29\] _04044_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout821_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10919__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06779_ _01905_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout919_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ _02165_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09498_ top.pc\[26\] _04518_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__or2_1
XANTENNA__07113__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08449_ _02495_ net488 net483 _02493_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _05288_ _05327_ _05287_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07416__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ net154 net2088 net329 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__mux2_1
XANTENNA__10654__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ top.a1.dataIn\[17\] _05257_ _05258_ top.a1.dataIn\[18\] _05259_ vssd1 vssd1
+ vccd1 vccd1 _05261_ sky130_fd_sc_hd__o221a_1
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13130_ clknet_leaf_37_clk _00694_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10342_ net1814 net247 net393 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13061_ clknet_leaf_118_clk _00625_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_52_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ net1587 net251 net403 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12012_ _05874_ _05881_ _05856_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__mux2_1
XANTENNA__07719__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13023__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout470 _03338_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_85_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12914_ clknet_leaf_51_clk _00478_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07352__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09892__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12845_ clknet_leaf_23_clk _00409_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_61_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10829__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ clknet_leaf_33_clk _00340_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08095__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06608__A _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ _05538_ _05575_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13865__1152 vssd1 vssd1 vccd1 vccd1 net1152 _13865__1152/LO sky130_fd_sc_hd__conb_1
XFILLER_0_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ _05526_ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ net147 net2113 net386 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10564__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ _05429_ _05455_ _05456_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold907 top.DUT.register\[13\]\[6\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__A2 _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold918 top.DUT.register\[22\]\[26\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ clknet_leaf_0_clk _00892_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold929 top.DUT.register\[10\]\[27\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_70_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06630__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13259_ clknet_leaf_29_clk _00823_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08907__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09654__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09580__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _02944_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__or2_4
XFILLER_0_209_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09580__B2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07591__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ net288 _02876_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ top.DUT.register\[24\]\[26\] net738 net717 top.DUT.register\[2\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a22o_1
XANTENNA__12746__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07682_ net809 _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__or2_1
XANTENNA__09883__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ _04459_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__nor2_1
X_06633_ top.DUT.register\[8\]\[28\] net569 net645 top.DUT.register\[17\]\[28\] _01759_
+ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a221o_1
XANTENNA_wire508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06697__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _04393_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__xnor2_1
X_06564_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ net481 net275 _03426_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09283_ _04328_ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__xnor2_1
X_06495_ top.a1.instruction\[31\] _01621_ net524 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__a21o_4
XFILLER_0_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ net276 _03251_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10982__B net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08165_ _03289_ _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__nor2_1
XANTENNA__10474__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout402_A _04939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07116_ top.DUT.register\[16\]\[12\] _01514_ _01539_ top.DUT.register\[13\]\[12\]
+ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08096_ _02731_ net289 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload80 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06621__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ top.DUT.register\[7\]\[10\] net684 net680 top.DUT.register\[13\]\[10\] _02173_
+ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a221o_1
Xclkload91 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout869_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A1 top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _03886_ _03902_ _03924_ _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_145_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09851__X _04850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _03054_ _03073_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_67_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ top.a1.row1\[61\] _04979_ _04986_ net849 vssd1 vssd1 vccd1 vccd1 _01118_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_3_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07334__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ top.pad.keyCode\[5\] top.pad.keyCode\[6\] top.pad.keyCode\[7\] top.pad.keyCode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__or4b_2
XANTENNA__06688__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10649__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net1573 net190 net348 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__mux2_1
X_12630_ clknet_leaf_2_clk _00194_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12561_ clknet_leaf_120_clk _00125_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _05381_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ clknet_leaf_99_clk _00059_ net982 vssd1 vssd1 vccd1 vccd1 top.ramstore\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11443_ _05246_ _05276_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10384__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06434__Y _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13275__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06163__A top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11374_ _05238_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and2_1
XANTENNA__08930__X _04026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_189_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ clknet_leaf_37_clk _00677_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10325_ top.DUT.register\[13\]\[22\] net184 net399 vssd1 vssd1 vccd1 vccd1 _00528_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_189_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06612__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ clknet_leaf_61_clk _00608_ net1099 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10256_ net1858 net184 net456 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__mux2_1
XANTENNA__11509__A top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10187_ net191 top.DUT.register\[9\]\[20\] net411 vssd1 vssd1 vccd1 vccd1 _00398_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07573__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11657__C1 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06679__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13877_ net1128 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12828_ clknet_leaf_55_clk _00392_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12759_ clknet_leaf_77_clk _00323_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06280_ net1469 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[24\] sky130_fd_sc_hd__and2_1
XFILLER_0_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09368__B top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06851__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06344__Y _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold704 top.DUT.register\[9\]\[25\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 top.DUT.register\[4\]\[30\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 top.DUT.register\[23\]\[31\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 top.DUT.register\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09970_ net1515 net237 net429 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
Xhold748 top.DUT.register\[17\]\[7\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06603__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold759 top.DUT.register\[22\]\[22\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ _03152_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__xnor2_1
XANTENNA_wire458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06360__X _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08852_ _03628_ _03770_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09671__X _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ top.DUT.register\[14\]\[19\] net614 net542 top.DUT.register\[22\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_108_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08783_ _01953_ _03884_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_127_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09305__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07734_ top.DUT.register\[25\]\[1\] net774 _01539_ top.DUT.register\[13\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11112__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10469__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ top.DUT.register\[8\]\[0\] net568 net623 top.DUT.register\[25\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout352_A _04963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _04446_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1094_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06616_ top.DUT.register\[25\]\[28\] net773 net741 top.DUT.register\[8\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a22o_1
X_07596_ top.DUT.register\[7\]\[3\] net681 net671 top.DUT.register\[16\]\[3\] _02722_
+ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _04380_ _04381_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06547_ top.DUT.register\[2\]\[30\] net660 net652 top.DUT.register\[28\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_173_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout617_A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ net823 _02210_ _02786_ _01615_ _01622_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__o221a_4
XANTENNA__07095__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06535__X _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ _01583_ net804 _01589_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08217_ net273 _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__or2_2
XFILLER_0_105_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ net908 top.pc\[7\] _04253_ net898 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09993__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _03272_ _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08595__A2 _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08079_ _01991_ net294 vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__or2_1
XANTENNA__10932__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08910__B net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10110_ net2341 net207 net462 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
X_11090_ net915 net1315 net853 _05031_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07085__Y _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ net226 net2280 net422 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__mux2_1
Xhold20 top.a1.hexop\[1\] vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _01176_ vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 top.a1.dataInTemp\[9\] vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top.lcd.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 top.a1.row1\[1\] vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold75 net100 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13800_ clknet_leaf_65_clk _01343_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold86 net124 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _01183_ vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11992_ _05836_ _05837_ _05846_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__nor3_1
XFILLER_0_203_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07307__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10943_ _01410_ _04973_ _04972_ _04970_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a211o_1
X_13731_ clknet_leaf_71_clk _01274_ net1093 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10874_ net1610 net253 net347 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_13662_ clknet_leaf_82_clk _01221_ net1011 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ clknet_leaf_118_clk _00177_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13593_ clknet_leaf_97_clk _01152_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09469__A _01929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12544_ clknet_leaf_80_clk _00108_ net1002 vssd1 vssd1 vccd1 vccd1 top.pc\[27\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07086__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06833__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[27\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[27\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__09188__B _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11426_ top.a1.dataIn\[17\] _05289_ _05290_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__and3_1
XANTENNA__09756__X _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11357_ _05223_ _05224_ _05201_ _05215_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__a211o_1
XANTENNA__10842__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ net1459 net247 net397 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
X_11288_ top.a1.row1\[12\] _05093_ _05097_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_169_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10414__Y _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ clknet_leaf_41_clk _00591_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ net1612 net246 net454 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__mux2_1
XANTENNA__06349__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07546__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1040 net1042 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
Xfanout1051 net1084 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07010__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1062 net1063 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1073 net1076 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 net39 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1095 net1097 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10289__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07450_ top.DUT.register\[29\]\[6\] net666 net658 top.DUT.register\[1\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XANTENNA__07171__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06401_ top.DUT.register\[25\]\[30\] net771 net721 top.DUT.register\[14\]\[30\] _01526_
+ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a221o_1
X_07381_ top.DUT.register\[2\]\[7\] net719 net675 top.DUT.register\[18\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09120_ _04169_ _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and2_1
X_06332_ _01332_ _01460_ _01333_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__and3b_1
XANTENNA__09379__A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08283__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ _03390_ _04067_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__nor2_1
X_06263_ net1415 net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[7\] sky130_fd_sc_hd__and2_1
XANTENNA__09098__B _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ top.DUT.register\[21\]\[31\] net574 net613 top.DUT.register\[14\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22o_1
XANTENNA__09666__X _04689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06194_ _01385_ _01411_ _01415_ _01419_ net1180 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
Xhold501 top.DUT.register\[22\]\[10\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 top.DUT.register\[12\]\[16\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 top.DUT.register\[7\]\[30\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold534 top.DUT.register\[13\]\[1\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 top.DUT.register\[5\]\[11\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10752__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold556 top.DUT.register\[25\]\[30\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06802__Y _01929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 top.DUT.register\[12\]\[24\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 top.DUT.register\[8\]\[28\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _04858_ net1797 net436 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__mux2_1
Xhold589 top.DUT.register\[24\]\[31\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
X_08904_ net276 _03961_ _04000_ _03201_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_5_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11149__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ net160 net2168 net437 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1107_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07001__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09842__A _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08835_ net474 _03924_ _03926_ net472 _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o221a_1
X_08766_ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__inv_2
X_07717_ top.DUT.register\[13\]\[1\] net649 net558 top.DUT.register\[6\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08697_ _03426_ _03542_ _03804_ net274 vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout734_A _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09988__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ top.DUT.register\[10\]\[2\] net727 _02772_ _02774_ vssd1 vssd1 vccd1 vccd1
+ _02775_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_49_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07579_ top.DUT.register\[8\]\[3\] net568 net619 top.DUT.register\[26\]\[3\] _02696_
+ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a221o_1
XANTENNA__10927__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ _04361_ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08265__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ net220 net1646 net387 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _04288_ _04289_ _04286_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_153_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ top.lcd.cnt_20ms\[9\] _06082_ net1107 vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ top.a1.row1\[13\] _05078_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__or2_1
X_12191_ _06049_ _06058_ _06050_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__o21a_1
XANTENNA__10662__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
X_11142_ net914 net1245 net854 _05057_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a31o_1
XANTENNA__07240__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06441__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_101_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__clkbuf_4
X_11073_ net89 net862 net826 net1188 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a22o_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__07528__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12431__RESET_B net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ net162 net2242 net425 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ _05840_ _05844_ _05828_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a21o_1
X_13714_ clknet_leaf_74_clk _01262_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ net177 net1805 net441 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ net1429 net194 net352 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XANTENNA__10837__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13645_ clknet_leaf_84_clk _01204_ net1014 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ net1526 net217 net445 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__mux2_1
X_13576_ clknet_leaf_96_clk _01135_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12527_ clknet_leaf_82_clk _00091_ net1013 vssd1 vssd1 vccd1 vccd1 top.pc\[10\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06806__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12458_ clknet_leaf_97_clk top.ru.next_FetchedInstr\[10\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ _05274_ _05277_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__xor2_1
XANTENNA__10572__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12389_ clknet_leaf_83_clk _00025_ net1014 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13317__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__RESET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06950_ _02056_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nor2_1
XANTENNA__07519__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ top.DUT.register\[4\]\[22\] net768 _01996_ _02007_ vssd1 vssd1 vccd1 vccd1
+ _02008_ sky130_fd_sc_hd__a211o_1
XANTENNA__08131__C_N _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08620_ net472 _03715_ _03717_ net475 _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__o221a_2
XANTENNA__09381__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08551_ _03664_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07502_ top.DUT.register\[8\]\[5\] net568 net540 top.DUT.register\[22\]\[5\] _02615_
+ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a221o_1
X_08482_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__inv_2
XANTENNA__11094__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09692__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13307__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07433_ top.DUT.register\[4\]\[6\] net768 net583 top.DUT.register\[12\]\[6\] _02559_
+ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a221o_1
XANTENNA__10747__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08725__B _03829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ _02485_ _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_102_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09103_ net534 _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06315_ _01456_ _01457_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07295_ _02418_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout315_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1057_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ _03999_ _04018_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06246_ net1635 net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[22\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_135_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07470__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09747__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold320 top.DUT.register\[12\]\[21\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10482__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold331 top.DUT.register\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ net1994 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
Xhold342 top.DUT.register\[12\]\[14\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 top.DUT.register\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 top.DUT.register\[7\]\[21\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold375 top.DUT.register\[21\]\[12\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout800 _04968_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_2
Xhold386 top.DUT.register\[12\]\[27\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 top.DUT.register\[13\]\[0\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _05025_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06430__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ net237 net2209 net433 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__mux2_1
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__buf_1
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_4
Xfanout844 _04966_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_2
Xfanout855 _01431_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09572__A _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_2
X_09867_ _04859_ _04862_ _01586_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 top.DUT.register\[23\]\[5\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_2
Xfanout899 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_2
XANTENNA_fanout949_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1031 top.DUT.register\[19\]\[30\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 top.pad.keyCode\[3\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net1342 net839 net817 _03919_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__a22o_1
Xhold1053 top.DUT.register\[12\]\[30\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08188__A _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1064 top.DUT.register\[24\]\[26\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _03813_ net340 net336 _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__o211a_2
XANTENNA__07930__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1075 top.DUT.register\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12834__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1086 top.DUT.register\[31\]\[29\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 top.DUT.register\[25\]\[12\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ _02037_ net470 _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _05578_ _05622_ _05623_ _05576_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a22o_1
XANTENNA__07289__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10711_ net252 net1681 net383 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _05556_ _05558_ _05557_ _05552_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__o211a_1
XANTENNA__10657__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13430_ clknet_leaf_119_clk _00994_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10642_ net141 net1872 net391 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06436__A _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ clknet_leaf_118_clk _00925_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08789__A2 _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ net167 net2066 net359 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07997__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net1381 _06113_ _06115_ net588 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__o211a_1
X_13292_ clknet_leaf_9_clk _00856_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09738__A1 _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ _06063_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__nor2_1
XANTENNA__10392__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07213__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12174_ _06019_ _06040_ _06042_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_75_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11125_ net54 net860 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ net102 net856 net825 net1267 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ net226 net1272 net428 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11236__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11958_ _05821_ _05823_ _05827_ _05819_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09674__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10284__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ net243 net1815 net443 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11889_ net129 _05749_ _05735_ _05740_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_15_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ clknet_leaf_61_clk net1228 net1101 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13559_ clknet_leaf_70_clk top.a1.nextHex\[2\] net1103 vssd1 vssd1 vccd1 vccd1 _01379_
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07988__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07080_ _02188_ _02205_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__or2_2
XANTENNA__07452__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06660__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08952__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout129 _05747_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
X_07982_ top.DUT.register\[9\]\[31\] net709 net706 top.DUT.register\[15\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09721_ net222 net2332 net439 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06933_ top.DUT.register\[11\]\[21\] net642 net606 top.DUT.register\[18\]\[21\] _02059_
+ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a221o_1
X_09652_ _01569_ net524 _01620_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__or3_4
X_06864_ _01982_ _01985_ _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__or3_4
XFILLER_0_179_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07912__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ _02361_ _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09583_ _01623_ net490 vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06795_ top.DUT.register\[19\]\[24\] net734 net669 top.DUT.register\[5\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ _03563_ _03648_ net304 vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08468__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ _03342_ _03582_ net312 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10477__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A _04920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ net809 _02540_ _02541_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ _02589_ _03515_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__nand2_1
XANTENNA__07691__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire508 _02254_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_162_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ top.DUT.register\[23\]\[8\] net560 net619 top.DUT.register\[26\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07443__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06543__X _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07278_ top.DUT.register\[4\]\[9\] net769 net683 top.DUT.register\[7\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09017_ _03584_ _03606_ _03626_ _03652_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout899_A top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06229_ net2353 net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[5\] sky130_fd_sc_hd__and2_1
XANTENNA__08190__B _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 _01197_ vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold161 top.ramstore\[27\] vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 top.ramaddr\[19\] vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 top.a1.row2\[3\] vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 top.ramstore\[2\] vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06403__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _01660_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_8
Xfanout641 _01648_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_8
X_09919_ _04909_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__xnor2_1
Xfanout652 _01641_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 _01636_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_8
Xfanout674 _01549_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 _01543_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_4
X_12930_ clknet_leaf_44_clk _00494_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout696 _01537_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07534__B _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ clknet_leaf_108_clk _00425_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11812_ _05672_ _05676_ top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_197_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12792_ clknet_leaf_107_clk _00356_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_194_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _05570_ _05611_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10387__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06166__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ _05492_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13413_ clknet_leaf_119_clk _00977_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06890__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10625_ net195 net1576 net391 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13344_ clknet_leaf_47_clk _00908_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ net233 net1292 net358 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06642__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10487_ net244 net2151 net368 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ clknet_leaf_53_clk _00839_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12226_ net1202 _06002_ net589 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_184_Right_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10850__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _06009_ _06023_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__xor2_2
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11108_ net914 net1271 net854 _05040_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a31o_1
X_12088_ _05896_ _05939_ _05932_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__mux2_1
X_11039_ net19 net842 net812 net1497 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06580_ top.DUT.register\[12\]\[29\] net582 _01699_ _01706_ vssd1 vssd1 vccd1 vccd1
+ _01707_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10297__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08250_ net313 _03374_ _03364_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07673__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__B2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07201_ top.DUT.register\[11\]\[15\] net756 net720 top.DUT.register\[14\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08181_ net503 net297 vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__nand2_1
XANTENNA__09658__Y _04681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07132_ top.DUT.register\[11\]\[12\] net641 net637 top.DUT.register\[16\]\[12\] _02258_
+ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07459__X _02586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07425__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08622__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08291__A _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06633__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07063_ net903 _01584_ _01609_ _02188_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10980__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10760__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _02037_ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout382_A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _02192_ _02204_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and2_1
X_06916_ top.DUT.register\[4\]\[21\] net768 net679 top.DUT.register\[13\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07896_ top.DUT.register\[6\]\[17\] net556 net623 top.DUT.register\[25\]\[17\] _03013_
+ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a221o_1
X_09635_ top.a1.halfData\[1\] _01472_ _04662_ net1103 vssd1 vssd1 vccd1 vccd1 _00117_
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ top.DUT.register\[6\]\[23\] net763 net716 top.DUT.register\[2\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ net138 _04585_ _04600_ net134 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o22a_1
X_06778_ net805 _01904_ _01624_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08466__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06538__X _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10248__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08517_ _02233_ _03612_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ _04527_ _04529_ _04526_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout814_A _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10000__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07664__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ net313 net482 _03565_ net469 _02496_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__o32a_1
XFILLER_0_147_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06872__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _03356_ _03360_ net306 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10410_ net156 net1798 net329 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__mux2_1
X_11390_ top.a1.dataIn\[18\] _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09381__A_N _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07416__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06624__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ net1917 net253 net394 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ clknet_leaf_39_clk _00624_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ net1663 net257 net402 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__mux2_1
X_12011_ _05874_ _05876_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_72_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10670__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_6
XFILLER_0_205_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_4
Xfanout482 _03184_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
X_12913_ clknet_leaf_12_clk _00477_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13893_ net1143 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_201_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12844_ clknet_leaf_10_clk _00408_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12775_ clknet_leaf_25_clk _00339_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11726_ _05534_ _05575_ _05537_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_83_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10845__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ _05500_ _05516_ _05520_ top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 _05527_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07407__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ net152 net2334 net388 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__mux2_1
X_11588_ _05455_ _05456_ _05429_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06615__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__C _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold908 top.DUT.register\[29\]\[28\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ clknet_leaf_23_clk _00891_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold919 top.DUT.register\[13\]\[20\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ net2306 net169 net363 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13258_ clknet_leaf_40_clk _00822_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13833__RESET_B net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__A2 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ top.a1.row2\[40\] net845 net813 _05750_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__a22o_1
XANTENNA__10580__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ clknet_leaf_120_clk _00753_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07040__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07750_ net288 _02876_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nor2_2
X_06701_ top.DUT.register\[6\]\[26\] net766 net698 top.DUT.register\[23\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a22o_1
X_07681_ _02804_ _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__or2_4
XFILLER_0_211_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06632_ top.DUT.register\[14\]\[28\] net613 net605 top.DUT.register\[18\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a22o_1
X_09420_ _04461_ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_189_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07894__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12786__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _04396_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__nor2_1
X_06563_ net806 _01689_ _01624_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08302_ net308 _03424_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__nand2_2
XFILLER_0_191_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ _04331_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__nor2_1
XANTENNA__08573__X _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06494_ _01477_ _01620_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__or2_2
XANTENNA__07646__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ net302 _03355_ _03357_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06854__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10755__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout228_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ _01713_ net293 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07115_ top.DUT.register\[12\]\[12\] net582 net698 top.DUT.register\[23\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a22o_1
X_08095_ net322 _03221_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload70 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__inv_8
XANTENNA__09845__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ top.DUT.register\[9\]\[10\] net711 net697 top.DUT.register\[23\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload81 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload92 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__inv_6
XANTENNA__08359__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10490__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06540__Y _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _03851_ _03867_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_145_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07948_ _03054_ _03073_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout931_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ top.DUT.register\[28\]\[17\] net584 _03004_ _03005_ vssd1 vssd1 vccd1 vccd1
+ _03006_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__B _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09618_ top.pad.keyCode\[1\] top.pad.keyCode\[0\] top.pad.keyCode\[3\] top.pad.keyCode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__or4b_2
XFILLER_0_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10890_ net1818 net193 net348 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ _04178_ _04574_ _04584_ _04044_ top.pc\[28\] vssd1 vssd1 vccd1 vccd1 _00109_
+ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_191_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08834__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07637__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ clknet_leaf_121_clk _00124_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08834__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11511_ _05379_ _05380_ _05375_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a21o_1
XANTENNA__10665__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_199_Left_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12491_ clknet_leaf_98_clk _00058_ net981 vssd1 vssd1 vccd1 vccd1 top.ramstore\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11442_ _05282_ _05310_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06444__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11373_ _05241_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_189_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10324_ net1787 net189 net399 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__mux2_1
X_13112_ clknet_leaf_109_clk _00676_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09755__A _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07270__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06731__X _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13043_ clknet_leaf_2_clk _00607_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10255_ net1479 net188 net456 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__mux2_1
XANTENNA__07022__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__A _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13350__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ net206 net1746 net410 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13876_ net1127 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__07876__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12827_ clknet_leaf_52_clk _00391_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07089__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ clknet_leaf_120_clk _00322_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06836__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ _05487_ _05529_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__or2_1
XANTENNA__10575__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12689_ clknet_leaf_12_clk _00253_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11188__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold705 top.DUT.register\[9\]\[14\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_203_Left_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold716 top.DUT.register\[11\]\[19\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 top.DUT.register\[11\]\[28\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09665__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold738 top.DUT.register\[30\]\[24\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07261__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold749 top.DUT.register\[3\]\[28\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ _01694_ _03997_ _01692_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__a21o_1
XANTENNA__07013__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08851_ _01820_ net486 net470 _01821_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a22o_1
XANTENNA__12598__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ top.DUT.register\[3\]\[19\] net788 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__and2_1
X_08782_ _01950_ _01951_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_127_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07733_ top.DUT.register\[17\]\[1\] net724 net718 top.DUT.register\[2\]\[1\] _02859_
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout178_A _04840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__A0 top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ top.DUT.register\[23\]\[0\] net560 net611 top.DUT.register\[14\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ _04422_ _04426_ _04427_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a21o_1
X_06615_ top.DUT.register\[4\]\[28\] net768 net586 top.DUT.register\[28\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__a22o_1
X_07595_ top.DUT.register\[14\]\[3\] net720 net716 top.DUT.register\[2\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout345_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ net136 _04372_ net907 vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__o21ai_1
X_06546_ top.DUT.register\[23\]\[30\] net561 net545 top.DUT.register\[5\]\[30\] _01672_
+ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a221o_1
XANTENNA__07619__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06827__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06477_ _01592_ _01593_ _01597_ _01603_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__and4_4
X_09265_ _04313_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10485__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08216_ net301 _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09196_ net137 _04243_ _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ _02099_ net293 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08078_ net514 net294 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__nand2_1
XANTENNA__13373__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ top.DUT.register\[7\]\[11\] net553 net783 top.DUT.register\[31\]\[11\] _02155_
+ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout979_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ net231 net1588 net422 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
XANTENNA__08201__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 top.a1.dataInTemp\[1\] vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 top.a1.dataInTemp\[6\] vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net115 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 top.ramstore\[0\] vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 net112 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _01172_ vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 top.ramaddr\[28\] vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__A _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 top.ramstore\[25\] vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ _05831_ _05857_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13730_ clknet_leaf_68_clk _01273_ vssd1 vssd1 vccd1 vccd1 top.lcd.lcd_rs sky130_fd_sc_hd__dfxtp_1
X_13879__1130 vssd1 vssd1 vccd1 vccd1 _13879__1130/HI net1130 sky130_fd_sc_hd__conb_1
X_10942_ net912 _01416_ _04967_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__or3b_1
XANTENNA__07858__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13661_ clknet_leaf_83_clk _01220_ net1017 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10873_ net1618 net255 net345 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ clknet_leaf_41_clk _00176_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13592_ clknet_leaf_96_clk _01151_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06818__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ clknet_leaf_89_clk _00107_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[26\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__10395__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07491__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ clknet_leaf_95_clk top.ru.next_FetchedInstr\[26\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _05289_ _05290_ top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08660__Y _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07243__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06461__X _01588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ _05223_ _05224_ _05215_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_111_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06597__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ net1996 net253 net399 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
X_11287_ net880 _05097_ _05098_ top.a1.row2\[12\] net879 vssd1 vssd1 vccd1 vccd1 _05163_
+ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_169_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ clknet_leaf_42_clk _00590_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ net2029 net251 net456 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_206_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_2
Xfanout1052 net1060 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
X_10169_ net259 net1782 net409 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
Xfanout1063 net1068 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1074 net1076 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_2
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09299__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13859_ net1150 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06400_ _01499_ net790 _01508_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__and3_4
XFILLER_0_186_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07380_ _02499_ _02501_ _02504_ _02506_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06331_ _01448_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06809__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ _03457_ _03485_ _03512_ _03534_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__and4_1
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06262_ top.ramload\[6\] net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_5_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08001_ top.DUT.register\[23\]\[31\] net562 net605 top.DUT.register\[18\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a22o_1
X_06193_ _01385_ _01415_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__nand2_1
XANTENNA__09223__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09223__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 top.DUT.register\[14\]\[20\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold513 top.DUT.register\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09395__A top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 top.DUT.register\[29\]\[25\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold535 top.DUT.register\[6\]\[4\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 top.DUT.register\[26\]\[26\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 top.DUT.register\[26\]\[4\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 top.DUT.register\[14\]\[18\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 top.DUT.register\[14\]\[11\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net173 net1982 net436 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__mux2_1
XANTENNA__06531__B net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08903_ _01713_ net291 net287 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _03955_ net343 _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_148_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08834_ net482 _03931_ _03932_ net519 _03934_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o221a_1
XANTENNA__09842__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1002_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ _03094_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06760__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07716_ top.DUT.register\[2\]\[1\] net662 net637 top.DUT.register\[16\]\[1\] _02842_
+ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__a221o_1
X_08696_ _03803_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07647_ top.DUT.register\[28\]\[2\] net584 net692 top.DUT.register\[21\]\[2\] _02773_
+ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_A _01523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07578_ _02697_ _02699_ _02701_ _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09317_ _04364_ _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06529_ _01573_ _01590_ net789 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__and3_2
XANTENNA__08265__A2 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07473__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _04298_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_153_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08017__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _04235_ _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ top.a1.state\[1\] _04978_ net530 net1283 vssd1 vssd1 vccd1 vccd1 _01263_
+ sky130_fd_sc_hd__a22o_1
X_12190_ _01399_ _06046_ _06052_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_186_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06579__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08973__B1 _01972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ net63 net858 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__and2_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
X_11072_ net1360 net856 net825 top.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 _01190_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XANTENNA__12889__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
X_10023_ net166 net2073 net427 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11088__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _05841_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__and2_1
XANTENNA__06169__A top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12400__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ clknet_leaf_74_clk _01261_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ net183 net1841 net443 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_127_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_197_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13644_ clknet_leaf_83_clk _01203_ net1017 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10856_ net1622 net204 net351 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13575_ clknet_leaf_96_clk _01134_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10787_ net1741 net227 net446 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__mux2_1
XANTENNA__07464__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ clknet_leaf_79_clk _00090_ net1004 vssd1 vssd1 vccd1 vccd1 top.pc\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ clknet_leaf_97_clk top.ru.next_FetchedInstr\[9\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[9\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10853__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08008__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11408_ _05274_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__nor2_1
XANTENNA__09756__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07216__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12388_ clknet_leaf_83_clk _00024_ net1017 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__B1 _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11339_ top.a1.dataIn\[22\] _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13009_ clknet_leaf_3_clk _00573_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06880_ top.DUT.register\[10\]\[22\] net729 net714 top.DUT.register\[30\]\[22\] _02002_
+ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a221o_1
XFILLER_0_206_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06742__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08550_ _02278_ _03663_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_145_Left_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07501_ _02619_ _02621_ _02623_ _02627_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__or4_1
X_08481_ _03373_ _03541_ _03585_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a211o_1
XANTENNA__09692__A1 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11713__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07432_ top.DUT.register\[6\]\[6\] net766 net717 top.DUT.register\[2\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07363_ _02486_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_170_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09102_ _02192_ _02198_ _02203_ _04152_ _02189_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__o41a_1
XANTENNA__07455__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06314_ _01333_ _01448_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07294_ top.DUT.register\[11\]\[9\] net756 net736 top.DUT.register\[24\]\[9\] _02415_
+ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a221o_1
XANTENNA__11251__B2 top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_198_Right_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08581__X _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06245_ top.ramload\[21\] net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09033_ _03715_ _03944_ _03992_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__and4_1
XFILLER_0_170_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10763__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Left_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07207__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06176_ net895 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
Xhold310 top.DUT.register\[13\]\[16\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12200__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 top.DUT.register\[13\]\[9\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 top.DUT.register\[11\]\[30\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 top.DUT.register\[24\]\[14\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 top.DUT.register\[12\]\[2\] vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__A0 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold365 top.DUT.register\[22\]\[7\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 top.DUT.register\[28\]\[27\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 top.DUT.register\[18\]\[7\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _01626_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_2
Xhold398 top.DUT.register\[14\]\[9\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout812 _05025_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_2
X_09935_ net239 net2187 net434 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__mux2_1
Xfanout823 _01565_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 _01567_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout677_A _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net847 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
Xfanout856 net861 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
Xfanout867 _01428_ vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_2
X_09866_ _04859_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_181_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 _01425_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_1
Xhold1010 top.DUT.register\[23\]\[14\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 top.DUT.register\[28\]\[28\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 net890 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_2
X_08817_ net889 top.pc\[25\] net537 _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a22o_1
Xhold1032 top.DUT.register\[30\]\[31\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1043 top.DUT.register\[4\]\[12\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 top.DUT.register\[12\]\[11\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _04797_ _04798_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__o21ai_2
Xhold1065 top.DUT.register\[22\]\[20\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 top.DUT.register\[5\]\[22\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09999__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1087 top.DUT.register\[24\]\[19\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _02036_ net487 net486 _02035_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a2bb2o_1
Xhold1098 top.DUT.register\[15\]\[16\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10817__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _03701_ _03787_ net304 vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__Y _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ net257 net1800 net381 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07694__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _01395_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ net144 net1537 net389 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06436__B _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07446__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ clknet_leaf_0_clk _00924_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_Left_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08643__C1 _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ net168 net2330 net360 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12311_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10673__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ clknet_leaf_29_clk _00855_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12242_ top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] top.lcd.cnt_20ms\[2\] vssd1 vssd1
+ vccd1 vccd1 _06073_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09738__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06452__A top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12173_ _06040_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_75_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11124_ net915 net1317 net853 _05048_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_166_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ net101 net862 net827 net1195 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_181_Left_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10006_ net234 net2309 net426 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06724__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10848__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11957_ _05817_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__and2b_1
XANTENNA__09674__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07685__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ net248 net1889 net441 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11888_ net129 _05749_ _05735_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__a21oi_2
X_13627_ clknet_leaf_45_clk net1270 net1081 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10839_ net1956 net259 net349 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_8__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_13558_ clknet_leaf_70_clk top.a1.nextHex\[1\] net1095 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08842__A _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ clknet_leaf_114_clk _00076_ net981 vssd1 vssd1 vccd1 vccd1 top.ramstore\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10583__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13489_ clknet_leaf_118_clk _01053_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08561__B _03483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07981_ top.DUT.register\[24\]\[31\] net737 net691 top.DUT.register\[3\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06963__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09720_ _03639_ net342 net336 _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__o211a_4
X_06932_ top.DUT.register\[25\]\[21\] net625 net598 top.DUT.register\[27\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a22o_1
XANTENNA__08289__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ top.pc\[1\] _04624_ _04674_ net897 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__o211a_1
X_06863_ _01987_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__or2_1
XANTENNA__06715__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ _02403_ _03691_ _02898_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a21oi_1
X_09582_ _01560_ _04606_ _04609_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__o21a_1
X_06794_ top.DUT.register\[30\]\[24\] net714 net676 top.DUT.register\[18\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
X_08533_ net277 _03602_ _03647_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10758__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout258_A _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _03477_ _03581_ net307 vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07140__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07415_ net809 _02540_ _02541_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_137_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _02589_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout425_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13181__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_2
X_07346_ top.DUT.register\[16\]\[8\] net635 net615 top.DUT.register\[30\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10493__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ _02320_ _02361_ _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__or3b_1
XANTENNA__08640__A2 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10983__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ _04023_ _04070_ _04071_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__or4_1
X_06228_ net1553 net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[4\] sky130_fd_sc_hd__and2_1
XFILLER_0_103_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08928__A0 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A _01492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 top.ramaddr\[0\] vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
X_06159_ top.edg2.flip2 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
Xhold151 top.DUT.register\[7\]\[28\] vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 top.DUT.register\[25\]\[11\] vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 top.ramload\[17\] vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 top.ramaddr\[1\] vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 top.DUT.register\[7\]\[20\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout961_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12801__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 _01663_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
XANTENNA__06954__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout631 _01656_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_4
Xfanout642 _01648_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_4
XANTENNA__11618__A top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ top.pc\[31\] _01623_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__xnor2_1
Xfanout653 _01641_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 _01636_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09870__X _04867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout675 _01549_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
Xfanout686 _01543_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
X_09849_ _04834_ _04837_ _04846_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_70_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout697 _01537_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ clknet_leaf_18_clk _00424_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07752__A_N _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ _05645_ _05677_ _05678_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a2bb2o_1
X_12791_ clknet_leaf_106_clk _00355_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10668__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07667__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ _05570_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06447__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07131__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11673_ _05465_ _05491_ _05466_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13412_ clknet_leaf_39_clk _00976_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07419__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ net200 net1938 net391 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13343_ clknet_leaf_115_clk _00907_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10555_ net235 net1840 net357 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13274_ clknet_leaf_19_clk _00838_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net247 net2027 net365 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12225_ net1297 _06018_ net589 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XANTENNA__07198__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _06024_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06945__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ net44 net858 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__and2_1
X_12087_ _05942_ _05947_ _05955_ _05941_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09780__X _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output54_A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ net18 net832 _05024_ net1469 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12420__Q top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_201_Right_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10578__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12989_ clknet_leaf_107_clk _00553_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06628__Y _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__B _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07460__B _02586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ top.DUT.register\[20\]\[15\] net747 net744 top.DUT.register\[31\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ _03304_ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07131_ top.DUT.register\[26\]\[12\] net621 net597 top.DUT.register\[27\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06363__Y _01492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06804__B net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07062_ _02188_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_132_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07830__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06397__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06936__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ _02080_ _03090_ _03087_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ _01613_ net342 net335 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a21boi_4
XANTENNA__08138__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ top.DUT.register\[28\]\[21\] net587 net733 top.DUT.register\[19\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a22o_1
X_07895_ top.DUT.register\[28\]\[17\] net651 net615 top.DUT.register\[30\]\[17\] _03021_
+ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_A _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _04650_ _04658_ _04659_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__or4_1
XANTENNA__07897__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ net805 _01972_ _01624_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a21o_1
XANTENNA__07361__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09565_ _04598_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10488__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout163_X net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ _01894_ _01903_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout542_A _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ _03629_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07649__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ _04532_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__or2_1
XANTENNA__08310__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07113__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08310__B2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08447_ _03544_ _03559_ _03558_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _03355_ _03366_ net298 vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07329_ top.DUT.register\[24\]\[8\] net735 net696 top.DUT.register\[23\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
XANTENNA__09271__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10340_ net1538 net256 net393 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07821__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10271_ net1514 net259 net401 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12010_ _05851_ _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_72_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 net453 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_6
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_6
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_4
XFILLER_0_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_2
X_12912_ clknet_leaf_122_clk _00476_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07888__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ net1142 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XANTENNA__07352__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ clknet_leaf_30_clk _00407_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10398__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06560__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11083__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_15__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ clknet_leaf_24_clk _00338_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11725_ _05581_ _05593_ _05574_ _05576_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_83_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08852__A2 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11656_ _05517_ _05518_ _05521_ _01394_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ net157 net1788 net387 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13326_ clknet_leaf_117_clk _00890_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold909 top.DUT.register\[21\]\[20\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ net1932 net172 net363 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07812__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13257_ clknet_leaf_2_clk _00821_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10861__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ net189 net2053 net371 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
XANTENNA__12997__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12208_ top.a1.row2\[35\] net845 net813 _05791_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__a22o_1
X_13188_ clknet_leaf_41_clk _00752_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06918__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _06007_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__or2_2
XANTENNA__07591__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06700_ top.DUT.register\[15\]\[26\] net707 _01535_ top.DUT.register\[3\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a22o_1
X_07680_ _02791_ _02792_ _02794_ _02806_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__or4_1
XFILLER_0_204_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08540__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08540__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ top.DUT.register\[15\]\[28\] _01655_ net783 top.DUT.register\[31\]\[28\]
+ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a221o_1
XANTENNA__06551__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ _03012_ _04394_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and2b_1
XANTENNA__10101__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06562_ _01673_ _01686_ _01687_ _01688_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__or4_4
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08301_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__inv_2
X_09281_ _02298_ _04329_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__and2b_1
XFILLER_0_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06493_ _01488_ net819 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__nand2_2
XFILLER_0_185_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08232_ net298 _03356_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11721__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08163_ _01560_ net297 vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__Y _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07114_ top.DUT.register\[28\]\[12\] net586 net702 top.DUT.register\[29\]\[12\] _02240_
+ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a221o_1
XANTENNA__07803__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08094_ _03204_ _03220_ net311 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload60 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10771__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07045_ top.DUT.register\[25\]\[10\] net771 net728 top.DUT.register\[10\]\[10\] _02169_
+ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a221o_1
Xclkload71 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload71/X sky130_fd_sc_hd__clkbuf_8
Xclkload82 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_6
XANTENNA__06821__Y _01948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ _03797_ _03819_ _03835_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06790__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A _01515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__Y _02779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ top.DUT.register\[26\]\[17\] net759 net674 top.DUT.register\[18\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a22o_1
XANTENNA__07334__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09617_ top.pad.keyCode\[5\] top.pad.keyCode\[4\] top.pad.keyCode\[7\] top.pad.keyCode\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__or4b_2
XANTENNA__11130__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06829_ top.DUT.register\[5\]\[23\] net544 net603 top.DUT.register\[18\]\[23\] _01955_
+ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout924_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09548_ net137 _04568_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__o22ai_1
XANTENNA__10011__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ top.a1.instruction\[25\] net822 _04424_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__o21a_2
XFILLER_0_136_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08834__A2 _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11510_ _05334_ _05376_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__xor2_2
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ clknet_leaf_62_clk _00057_ net1101 vssd1 vssd1 vccd1 vccd1 top.ramstore\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07320__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12496__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06444__B _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ _05209_ _05230_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13111_ clknet_leaf_77_clk _00675_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10323_ net2079 net193 net399 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10681__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__B1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ clknet_leaf_50_clk _00606_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ net1399 net191 net457 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__mux2_1
X_10185_ net214 net1566 net411 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
XANTENNA__07573__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
XANTENNA__08658__Y _03768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout291 net293 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06459__X _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07325__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__RESET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13875_ net1126 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_158_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12826_ clknet_leaf_19_clk _00390_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12757_ clknet_leaf_8_clk _00321_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10856__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__Y _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ clknet_leaf_122_clk _00252_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _05504_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 top.DUT.register\[4\]\[24\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 top.DUT.register\[14\]\[7\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_108_clk _00873_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold728 top.DUT.register\[17\]\[15\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10591__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold739 top.DUT.register\[10\]\[9\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
X_08850_ net314 net284 _03410_ _03545_ _03745_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o311a_1
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08849__X _03949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ _02921_ _02927_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__nor2_8
X_08781_ _01992_ _03866_ _01993_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06772__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07732_ top.DUT.register\[14\]\[1\] net723 net669 top.DUT.register\[5\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XANTENNA__08513__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11112__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08513__B2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09710__B1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07663_ top.DUT.register\[5\]\[0\] net544 net540 top.DUT.register\[22\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ _04444_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_140_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06614_ top.DUT.register\[21\]\[28\] net694 net687 top.DUT.register\[1\]\[28\] _01740_
+ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07594_ top.DUT.register\[12\]\[3\] net580 net726 top.DUT.register\[17\]\[3\] _02713_
+ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a221o_1
X_09333_ _04361_ _04365_ _04363_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06545_ top.DUT.register\[16\]\[30\] net636 net541 top.DUT.register\[22\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10766__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09264_ _04314_ _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06476_ _01598_ _01599_ _01600_ _01602_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ net286 _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ net133 _04248_ _04250_ _04251_ net908 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__o221a_1
X_08146_ _02810_ _02928_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08077_ net302 _03203_ _03198_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07028_ top.DUT.register\[19\]\[11\] net633 _01682_ top.DUT.register\[15\]\[11\]
+ _02144_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a221o_1
XFILLER_0_178_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 top.a1.dataInTemp\[2\] vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 net110 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 top.a1.row1\[9\] vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net1329 net868 _01731_ net594 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 top.a1.row1\[0\] vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 _01167_ vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06763__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 top.a1.dataInTemp\[7\] vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold77 top.a1.row1\[10\] vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 top.lcd.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ top.a1.dataIn\[4\] _05848_ _05859_ _05851_ vssd1 vssd1 vccd1 vccd1 _05860_
+ sky130_fd_sc_hd__or4b_4
Xhold99 _01192_ vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ net851 _04971_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__nor2_1
XANTENNA__08000__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_203_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660_ clknet_leaf_83_clk _01219_ net1011 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ net1820 net260 net345 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12611_ clknet_leaf_41_clk _00175_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_117_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13591_ clknet_leaf_97_clk _01150_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10676__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ clknet_leaf_102_clk _00106_ net1002 vssd1 vssd1 vccd1 vccd1 top.pc\[25\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_19_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[25\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11424_ _05292_ _05293_ _05260_ _05291_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09768__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09244__A_N _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11355_ _05223_ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10306_ net1869 net258 net400 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11286_ net880 _05097_ net879 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13465__RESET_B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ clknet_leaf_27_clk _00589_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ net1305 net255 net454 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__mux2_1
Xfanout1020 net39 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_2
XANTENNA__09940__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07546__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1031 net1038 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1051 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_2
Xfanout1053 net1060 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_58_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10168_ net264 net1591 net410 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XANTENNA__06754__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1067 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1086 net1110 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_2
Xfanout1097 net1110 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_2
X_10099_ net1425 net264 net461 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_179_Right_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13858_ net1149 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_186_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08845__A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12809_ clknet_leaf_4_clk _00373_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_108_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13789_ clknet_leaf_67_clk _01332_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_06330_ _01447_ _01468_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06261_ net2353 net878 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[5\] sky130_fd_sc_hd__and2_1
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ net490 vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__inv_2
X_06192_ net1401 _01419_ _01420_ top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 _00009_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold503 top.DUT.register\[12\]\[3\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09395__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 top.a1.row2\[2\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold525 top.DUT.register\[27\]\[18\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold536 top.DUT.register\[2\]\[26\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 top.ramload\[14\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold558 top.DUT.register\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ net177 net2137 net433 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
Xhold569 top.DUT.register\[9\]\[23\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ _01694_ _03105_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__xor2_1
XANTENNA__10902__X _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _04875_ _04876_ _04877_ net339 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_5_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07537__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ _01863_ net488 _03607_ _03771_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout190_A _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08764_ _01994_ _03093_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__or2_1
X_07715_ top.DUT.register\[7\]\[1\] net554 net597 top.DUT.register\[27\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__a22o_1
X_08695_ _03724_ _03802_ net307 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout455_A _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07646_ top.DUT.register\[4\]\[2\] net767 net755 top.DUT.register\[11\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10496__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ top.DUT.register\[21\]\[3\] net572 net599 top.DUT.register\[10\]\[3\] _02703_
+ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout622_A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ _02339_ _04362_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__and2b_1
X_06528_ net900 _01590_ _01591_ net801 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__and4b_4
XFILLER_0_192_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06275__A top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ top.pc\[10\] _02428_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06459_ net904 net823 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12199__A2_N _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ _04218_ _04221_ _04219_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06562__X _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08490__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08129_ net479 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12216__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_186_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140_ net914 net1331 net854 _05056_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__a31o_1
XANTENNA__06984__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XANTENNA__06733__A_N _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
X_11071_ net87 net862 net826 net1222 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a22o_1
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07528__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ net170 net1511 net426 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _05813_ _05838_ _05842_ _05805_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ net189 net1879 net443 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
X_13712_ clknet_leaf_73_clk _01260_ net1091 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07161__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07700__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10855_ net2025 net211 net352 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
X_13643_ clknet_leaf_86_clk _01202_ net1007 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11091__A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11245__C1 _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13574_ clknet_leaf_96_clk _01133_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ top.DUT.register\[27\]\[15\] net179 net445 vssd1 vssd1 vccd1 vccd1 _00969_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12525_ clknet_leaf_79_clk _00089_ net1004 vssd1 vssd1 vccd1 vccd1 top.pc\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12456_ clknet_leaf_100_clk top.ru.next_FetchedInstr\[8\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _05244_ _05245_ _05246_ _05256_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or4b_2
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12387_ clknet_leaf_83_clk _00023_ net1014 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11338_ _05189_ _05193_ top.a1.dataIn\[21\] top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 _05208_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_50_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08964__B2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__Q top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ net1246 net824 _05146_ net1090 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08399__X _03520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07519__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ clknet_leaf_0_clk _00572_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06727__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07500_ top.DUT.register\[29\]\[5\] net663 _02625_ _02626_ vssd1 vssd1 vccd1 vccd1
+ _02627_ sky130_fd_sc_hd__a211o_1
XANTENNA__07750__Y _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _03367_ net270 net268 _03358_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12528__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__A _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__A2 _01492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07431_ top.DUT.register\[8\]\[6\] net742 _02548_ _02557_ vssd1 vssd1 vccd1 vccd1
+ _02558_ sky130_fd_sc_hd__a211o_1
XANTENNA__11713__B top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06606__A_N _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07362_ top.DUT.register\[24\]\[8\] net548 net544 top.DUT.register\[5\]\[8\] _02474_
+ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ _04155_ _04158_ _04161_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__a21o_1
X_06313_ _01453_ _01455_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07293_ top.DUT.register\[13\]\[9\] net680 net668 top.DUT.register\[5\]\[9\] _02419_
+ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09032_ _03870_ _03972_ _04092_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__and4_1
X_06244_ net2156 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[20\] sky130_fd_sc_hd__and2_1
XANTENNA__06382__X _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06823__A _01929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 top.DUT.register\[1\]\[14\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06175_ top.Wen vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
Xhold311 top.DUT.register\[14\]\[19\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 top.DUT.register\[9\]\[13\] vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold333 top.ramaddr\[12\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold344 top.DUT.register\[27\]\[8\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold355 top.DUT.register\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 top.DUT.register\[27\]\[17\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 top.DUT.register\[22\]\[30\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout802 net804 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_2
Xhold388 top.DUT.register\[25\]\[16\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 top.DUT.register\[8\]\[22\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net243 net1874 net435 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__mux2_1
XANTENNA__09853__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06430__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout813 _04975_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
Xfanout824 _01443_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
Xfanout835 _01567_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09904__B1 _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07654__A _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net861 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_2
X_09865_ _04860_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__nand2_1
XANTENNA__06718__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 top.DUT.register\[4\]\[3\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_181_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout572_A _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_2
Xhold1011 top.DUT.register\[18\]\[29\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 top.pad.keyCode\[0\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 top.DUT.register\[19\]\[6\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _03916_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__nand2_1
Xhold1044 top.DUT.register\[20\]\[11\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ net834 _04415_ _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__o21ba_1
Xhold1055 top.DUT.register\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 top.DUT.register\[22\]\[8\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ net314 _03498_ _03745_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__o21ai_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 top.DUT.register\[31\]\[3\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 top.DUT.register\[7\]\[2\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08678_ _03746_ _03786_ net278 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07629_ top.DUT.register\[20\]\[2\] net576 net647 top.DUT.register\[13\]\[2\] _02744_
+ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10640_ net153 net1835 net391 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08643__B1 _03742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ net173 net1554 net358 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12310_ _01439_ _06109_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07997__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ clknet_leaf_34_clk _00854_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ _06071_ _06072_ net1108 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12172_ _06034_ _06035_ _06036_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11123_ net53 net859 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07564__A _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ net1235 net856 net825 top.ramstore\[5\] vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__a22o_1
X_10005_ net235 net2312 net425 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07382__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08666__Y _03776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11956_ _05822_ _05823_ _05815_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a21boi_1
XANTENNA__07134__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__A _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09674__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06908__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ net252 net2045 net443 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11887_ _05755_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ clknet_leaf_61_clk net1240 net1101 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10838_ net1406 net265 net351 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12418__Q top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13557_ clknet_leaf_69_clk top.a1.nextHex\[0\] net1103 vssd1 vssd1 vccd1 vccd1 _01378_
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10864__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ net146 net2085 net374 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07988__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ clknet_leaf_61_clk _00075_ net1099 vssd1 vssd1 vccd1 vccd1 top.ramstore\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13488_ clknet_leaf_0_clk _01052_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ clknet_leaf_94_clk top.ru.next_FetchedData\[23\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12194__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _01560_ _01691_ _03106_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_130_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06931_ top.DUT.register\[10\]\[21\] net601 net543 top.DUT.register\[22\]\[21\] _02057_
+ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08289__B _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09650_ _04045_ _04186_ _04671_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a31o_1
XANTENNA__10104__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ top.DUT.register\[24\]\[23\] net735 net726 top.DUT.register\[17\]\[23\] _01988_
+ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a221o_1
XANTENNA__07373__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ net1555 net839 net815 _03713_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a22o_1
XANTENNA__07912__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ net908 top.pc\[30\] _04610_ _04614_ net897 vssd1 vssd1 vccd1 vccd1 _00111_
+ sky130_fd_sc_hd__o221a_1
X_06793_ top.DUT.register\[25\]\[24\] net774 net718 top.DUT.register\[2\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
X_08532_ net287 _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06377__X _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08509__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07125__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08965__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _03535_ _03580_ net281 vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ net809 _02521_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nand2_1
X_08394_ _03450_ _03514_ _02634_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_137_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10432__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08244__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ _02400_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _04004_ _03985_ _03968_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06227_ net1359 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[3\] sky130_fd_sc_hd__and2_1
XANTENNA__08928__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ net901 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
Xhold141 top.ramaddr\[3\] vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 top.ramaddr\[20\] vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 top.DUT.register\[7\]\[13\] vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 top.a1.row1\[122\] vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06403__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold185 top.a1.row2\[11\] vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__B net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 top.pad.button_control.r_counter\[14\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _01667_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_4
Xfanout621 _01663_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_8
Xfanout632 _01656_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_2
X_09917_ top.pc\[30\] _04605_ _04903_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__a21o_1
Xfanout643 _01647_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_4
Xfanout654 _01641_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09353__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 _01636_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_8
Xfanout676 _01549_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10014__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09848_ _04834_ _04837_ _04846_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a21o_1
Xfanout687 _01543_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout698 _01537_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ net335 _04782_ _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_161_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A1 _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11810_ top.a1.dataIn\[7\] _05619_ _05642_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or3b_1
X_12790_ clknet_leaf_120_clk _00354_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07116__B1 _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11741_ _05549_ _05572_ _05599_ _05601_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__o31a_1
XFILLER_0_178_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06447__B top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11672_ _05516_ _05521_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09408__A2 top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10623_ net208 net2315 net391 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__mux2_1
X_13411_ clknet_leaf_22_clk _00975_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10684__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06890__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13342_ clknet_leaf_14_clk _00906_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10554_ net239 net2262 net360 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__A1 top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__B2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ clknet_leaf_36_clk _00837_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06642__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10485_ net251 net1643 net367 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__mux2_1
XANTENNA__06182__B _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ net1226 _06028_ net589 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
X_12155_ _06004_ _06009_ _06016_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__nor3_1
XFILLER_0_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ net917 net1493 net852 _05039_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a31o_1
X_12086_ _05942_ _05947_ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_88_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11037_ net17 net841 net811 net1424 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__o22a_1
XANTENNA__07355__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09713__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10859__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12988_ clknet_leaf_55_clk _00552_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11939_ _05775_ _05786_ _05790_ _05767_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13609_ clknet_leaf_61_clk net1265 net1100 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10594__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06881__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_12_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07130_ top.DUT.register\[8\]\[12\] net569 net644 top.DUT.register\[17\]\[12\] _02256_
+ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07061_ _01596_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__nor2_1
XANTENNA__06633__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07594__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _02122_ _03086_ _03088_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_79_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06914_ top.DUT.register\[2\]\[21\] net717 net691 top.DUT.register\[3\]\[21\] _02040_
+ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ top.a1.dataIn\[7\] _04716_ net343 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a21o_1
X_07894_ top.DUT.register\[2\]\[17\] net659 net619 top.DUT.register\[26\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a22o_1
XANTENNA__12543__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07346__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ _04643_ _04653_ _04648_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a21oi_1
X_06845_ _01956_ _01969_ _01970_ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__or4_4
XANTENNA__10769__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A _04959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _04569_ _04570_ _04571_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__o21ai_1
X_06776_ _01896_ _01898_ _01900_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_143_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08515_ net284 _03410_ _03544_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09495_ top.pc\[26\] _04515_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08310__A2 _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ _03186_ _03564_ net310 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__mux2_2
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06872__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08377_ _03494_ _03497_ net283 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__mux2_1
XANTENNA__09578__B _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07328_ top.DUT.register\[6\]\[8\] net763 net681 top.DUT.register\[7\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12649__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06624__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07259_ top.DUT.register\[23\]\[14\] net563 net542 top.DUT.register\[22\]\[14\] _02385_
+ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a221o_1
XANTENNA__07821__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10009__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ net1582 net264 net403 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout440 _04681_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
Xfanout451 net453 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_21_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout462 _04928_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_4
Xfanout473 _03335_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_4
XANTENNA__07337__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout484 _03180_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_2
X_12911_ clknet_leaf_22_clk _00475_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10679__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891_ net1141 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_88_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12842_ clknet_leaf_34_clk _00406_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06458__A top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12773_ clknet_leaf_116_clk _00337_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13424__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11724_ _05581_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11655_ _05446_ _05488_ _05523_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10606_ net162 net1948 net385 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__mux2_1
X_11586_ _05395_ _05426_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__xor2_2
XANTENNA__06615__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537_ net1420 net177 net361 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13325_ clknet_leaf_23_clk _00889_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10468_ net193 net1595 net372 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__mux2_1
X_13256_ clknet_leaf_33_clk _00820_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ top.a1.row2\[34\] net845 net813 _05824_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__a22o_1
X_13187_ clknet_leaf_41_clk _00751_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10399_ net217 net2233 net327 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__mux2_1
XANTENNA__07576__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09009__A _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ _05981_ _05993_ _06002_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__and3_1
XANTENNA__07040__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12431__Q top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ _05908_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_193_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07328__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06630_ top.DUT.register\[19\]\[28\] net633 net787 top.DUT.register\[3\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06368__A _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire503_A _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06561_ top.DUT.register\[8\]\[30\] net571 net600 top.DUT.register\[10\]\[30\] _01674_
+ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ net281 _03340_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09280_ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06492_ top.a1.instruction\[2\] _01494_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nand2_4
XFILLER_0_129_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08231_ _03244_ _03248_ net279 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06854__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08162_ _03287_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07113_ top.DUT.register\[20\]\[12\] net749 net730 top.DUT.register\[10\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ _03219_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_12
X_07044_ top.DUT.register\[12\]\[10\] net580 net726 top.DUT.register\[17\]\[10\] _02170_
+ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a221o_1
XANTENNA__06390__X _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload61 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload72 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_8
XANTENNA__12795__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload83 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload94 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_8
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12724__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ _03760_ _03782_ _04056_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout485_A _03179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07946_ net807 _03072_ _01624_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_145_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07662__A _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ top.DUT.register\[10\]\[17\] net727 net708 top.DUT.register\[9\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout652_A _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ top.pad.keyCode\[1\] top.pad.keyCode\[2\] top.pad.keyCode\[3\] top.pad.keyCode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_3_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06828_ top.DUT.register\[16\]\[23\] net635 net627 top.DUT.register\[9\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ _04575_ _04581_ _01618_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o21ai_1
X_06759_ top.DUT.register\[20\]\[25\] net577 net616 top.DUT.register\[30\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout917_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10626__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _04515_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08429_ _02587_ _03516_ _03525_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload0 clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
X_11440_ _05289_ _05290_ _05272_ _05280_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_156_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__A1 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11371_ _05203_ _05240_ _05239_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13110_ clknet_leaf_121_clk _00674_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10322_ net1371 net205 net398 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_189_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13041_ clknet_leaf_110_clk _00605_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ net1876 net205 net455 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__mux2_1
XANTENNA__07556__B _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06460__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ net215 net2271 net409 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_208_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07843__Y _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11106__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 _03238_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_4
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_2
XFILLER_0_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10202__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13874_ top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ clknet_leaf_37_clk _00389_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07089__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ clknet_leaf_60_clk _00320_ net1102 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ _05574_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06836__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12687_ clknet_leaf_21_clk _00251_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11638_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12426__Q top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10872__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11569_ _05404_ _05437_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 top.DUT.register\[15\]\[26\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_53_clk _00872_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold718 top.a1.row1\[111\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 top.DUT.register\[31\]\[5\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07261__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13239_ clknet_leaf_17_clk _00803_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07013__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__C_N _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _02911_ _02912_ _02924_ _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__or4_4
X_08780_ net1166 net840 net815 _03883_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07482__A top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07731_ top.DUT.register\[15\]\[1\] net706 net695 top.DUT.register\[21\]\[1\] _02857_
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07662_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__inv_2
XANTENNA__09710__B2 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06524__A1 top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06613_ top.DUT.register\[10\]\[28\] net729 net673 top.DUT.register\[16\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ _04443_ net512 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_140_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07593_ top.DUT.register\[8\]\[3\] net739 net700 top.DUT.register\[29\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06544_ _01628_ net789 _01637_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__and3_4
X_09332_ _03054_ _04378_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09263_ net894 _04304_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_173_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06475_ _01561_ _01601_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__nor2_1
XANTENNA__06827__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13720__Q top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08214_ _02831_ _03316_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ _04233_ _04237_ _04249_ _01619_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08145_ _03267_ _03270_ net282 vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10782__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ _03200_ _03202_ net288 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09529__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07027_ top.DUT.register\[11\]\[11\] net642 net609 top.DUT.register\[12\]\[11\] _02145_
+ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08201__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07004__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 top.pad.button_control.r_counter\[16\] vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 top.ramstore\[8\] vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net518 net592 net1198 net869 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__a2bb2o_1
Xhold34 net114 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 top.a1.row1\[19\] vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 net113 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 top.ramstore\[20\] vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 top.a1.dataInTemp\[10\] vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ top.DUT.register\[7\]\[16\] net555 net624 top.DUT.register\[25\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__a22o_1
Xhold89 top.lcd.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10022__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ top.a1.state\[2\] top.a1.state\[0\] top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04971_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08775__X _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ net1413 net263 net347 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12610_ clknet_leaf_42_clk _00174_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06295__X _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ clknet_leaf_98_clk _01149_ net982 vssd1 vssd1 vccd1 vccd1 top.ramload\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06736__A _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ clknet_leaf_102_clk _00105_ net997 vssd1 vssd1 vccd1 vccd1 top.pc\[24\] sky130_fd_sc_hd__dfstp_2
XANTENNA__06818__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6__f_clk_X clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[24\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[24\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07491__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09768__A1 _03757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11423_ top.a1.dataIn\[17\] _05235_ _05257_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__or3_1
XANTENNA__10692__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11354_ top.a1.dataIn\[31\] _05194_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__nand2_4
XANTENNA__06471__A top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07243__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10305_ net1752 net260 net397 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XANTENNA__11089__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ _05105_ _05116_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__or2_1
X_13024_ clknet_leaf_49_clk _00588_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10236_ net1837 net260 net454 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__mux2_1
XANTENNA__09782__A top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1010 net1012 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
X_10167_ net148 top.DUT.register\[9\]\[0\] net409 vssd1 vssd1 vccd1 vccd1 _00378_
+ sky130_fd_sc_hd__mux2_1
Xfanout1032 net1038 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08398__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1065 net1067 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_4
Xfanout1076 net1084 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_2
XFILLER_0_89_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10098_ net2291 net151 net459 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1087 net1110 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_4
Xfanout1098 net1109 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09006__B _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09721__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13857_ net1148 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_202_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10867__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12808_ clknet_leaf_32_clk _00372_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13788_ clknet_leaf_67_clk _01331_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06809__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12739_ clknet_leaf_50_clk _00303_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06260_ net1553 net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[4\] sky130_fd_sc_hd__and2_1
XFILLER_0_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13142__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06191_ _01413_ _01419_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nor2_1
XANTENNA__07748__Y _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold504 top.DUT.register\[30\]\[11\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold515 top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08431__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06381__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold526 top.DUT.register\[27\]\[29\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold537 top.DUT.register\[13\]\[29\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 top.DUT.register\[27\]\[7\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09950_ net186 net1971 net435 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__mux2_1
Xhold559 top.DUT.register\[12\]\[26\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10107__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08901_ _01694_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__xnor2_1
X_09881_ _04557_ net526 net332 top.a1.dataIn\[27\] net334 vssd1 vssd1 vccd1 vccd1
+ _04877_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08579__Y _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08832_ _01865_ _03338_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__nand2_1
XANTENNA__07942__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__C _03844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ _01994_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08101__A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13175__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ top.DUT.register\[20\]\[1\] net578 net569 top.DUT.register\[8\]\[1\] _02840_
+ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a221o_1
X_08694_ _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__inv_2
XANTENNA__08498__B2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10777__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ top.DUT.register\[30\]\[2\] net712 net671 top.DUT.register\[16\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout350_A _04963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ top.DUT.register\[1\]\[3\] net655 net781 top.DUT.register\[31\]\[3\] _02702_
+ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06527_ _01590_ _01628_ _01631_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__and3_1
X_09315_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout615_A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06458_ top.a1.instruction\[5\] _01565_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__nor2_1
X_09246_ top.pc\[10\] _02428_ _04283_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07473__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06681__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _04233_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nand2_1
X_06389_ _01499_ net792 _01506_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08128_ _03164_ _03182_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08059_ net300 _03185_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_186_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10017__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
X_11070_ net1284 net862 net826 top.ramstore\[21\] vssd1 vssd1 vccd1 vccd1 _01188_
+ sky130_fd_sc_hd__a22o_1
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XANTENNA__07460__A_N _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__08489__Y _03606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net174 net1866 net426 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
XANTENNA__09922__A1 top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ _05822_ _05823_ _05802_ _05808_ _05812_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11088__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_73_clk _01259_ net1093 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10923_ net191 net1950 net444 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10687__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13642_ clknet_leaf_83_clk _01201_ net1011 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
X_10854_ net2183 net216 net349 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
XANTENNA__09438__B1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06466__A top.a1.instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ clknet_leaf_85_clk _01132_ net1018 vssd1 vssd1 vccd1 vccd1 top.a1.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06185__B top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10785_ net1407 net196 net447 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09777__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12524_ clknet_leaf_78_clk _00088_ net1004 vssd1 vssd1 vccd1 vccd1 top.pc\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_137_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07464__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06672__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ clknet_leaf_100_clk top.ru.next_FetchedInstr\[7\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ _05245_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__or2_1
XANTENNA__08413__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07216__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ clknet_leaf_82_clk _00022_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06424__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11337_ _05204_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07584__X _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ _05139_ _05141_ _05143_ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__or4_1
XANTENNA__09913__A1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ clknet_leaf_22_clk _00571_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10219_ net213 top.DUT.register\[10\]\[18\] net408 vssd1 vssd1 vccd1 vccd1 _00428_
+ sky130_fd_sc_hd__mux2_1
X_11199_ net850 _05073_ net531 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__and3_1
XANTENNA__07924__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07953__A_N _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09017__A _03584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09677__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10597__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07430_ top.DUT.register\[9\]\[6\] net710 net682 top.DUT.register\[7\]\[6\] _02556_
+ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11713__C top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07361_ top.DUT.register\[6\]\[8\] net556 net540 top.DUT.register\[22\]\[8\] _02487_
+ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06312_ _01332_ _01452_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__or2_1
X_09100_ _04155_ _04158_ _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_102_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07455__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07292_ top.DUT.register\[25\]\[9\] net771 net740 top.DUT.register\[8\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ _03671_ _03692_ _03846_ _03863_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__and4_1
X_06243_ top.ramload\[19\] net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[19\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06174_ top.Ren vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XANTENNA__07207__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12200__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 top.DUT.register\[29\]\[31\] vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 top.a1.hexop\[4\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 top.DUT.register\[11\]\[23\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06415__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold334 top.DUT.register\[14\]\[1\] vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 top.DUT.register\[23\]\[12\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 top.DUT.register\[19\]\[15\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top.DUT.register\[13\]\[14\] vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 top.DUT.register\[14\]\[3\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net248 net2272 net433 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__mux2_1
Xhold389 top.DUT.register\[30\]\[15\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout814 _04975_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_209_Left_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13038__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout825 net829 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_2
XANTENNA__09904__A1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 _01567_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07654__B _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ top.pc\[26\] _04543_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__or2_1
Xfanout847 _04635_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
Xfanout858 net860 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_2
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_181_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 top.DUT.register\[15\]\[18\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1105_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 top.DUT.register\[21\]\[13\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _03898_ _03915_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1023 top.DUT.register\[29\]\[17\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _04425_ net526 net333 top.a1.dataIn\[19\] net334 vssd1 vssd1 vccd1 vccd1
+ _04799_ sky130_fd_sc_hd__a221o_1
Xhold1034 top.DUT.register\[13\]\[15\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 top.DUT.register\[8\]\[20\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 top.DUT.register\[24\]\[2\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 top.DUT.register\[18\]\[20\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ _02037_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09668__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1078 top.a1.data\[3\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 top.DUT.register\[16\]\[30\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
X_08677_ _03212_ _03216_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08340__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ top.DUT.register\[24\]\[2\] net548 net603 top.DUT.register\[18\]\[2\] _02745_
+ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__a221o_1
XANTENNA__10300__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07694__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12991__RESET_B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ top.a1.instruction\[10\] _01477_ _01620_ top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _02686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10570_ net175 net2117 net357 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__mux2_1
XANTENNA__07446__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08643__A1 _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08643__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06654__B1 _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ top.pc\[9\] _02472_ _04276_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06733__B _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _06072_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_161_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12171_ _06031_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_75_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ net916 net1312 net854 _05047_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a31o_1
Xhold890 top.DUT.register\[12\]\[28\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11053_ net99 net864 net828 net1274 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ net241 net2256 net425 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
XANTENNA__08947__Y _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11955_ _05792_ _05823_ _05821_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__mux2_2
XANTENNA__06908__B _02034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ net258 net2237 net441 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XANTENNA__10210__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07685__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ _05702_ _05738_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06893__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ clknet_leaf_114_clk net1261 net940 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
X_10837_ net2147 net149 net349 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ clknet_leaf_72_clk _01120_ net1104 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[63\]
+ sky130_fd_sc_hd__dfstp_1
X_10768_ net152 net2325 net375 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09300__A _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06645__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12507_ clknet_leaf_100_clk _00074_ net986 vssd1 vssd1 vccd1 vccd1 top.ramstore\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13487_ clknet_leaf_20_clk _01051_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ net174 net1628 net378 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12438_ clknet_leaf_94_clk top.ru.next_FetchedData\[22\] net995 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10880__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ net795 _06150_ _06151_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09347__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ top.DUT.register\[2\]\[21\] net661 net613 top.DUT.register\[14\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a22o_1
X_06861_ top.DUT.register\[27\]\[23\] net775 net712 top.DUT.register\[30\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a22o_1
XANTENNA__08570__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ net886 top.pc\[14\] net539 _03712_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__a22o_1
X_09580_ net138 _04604_ _04613_ net133 net908 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o221ai_1
X_06792_ _01913_ _01915_ _01917_ _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__or4_2
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08531_ _03242_ _03247_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08322__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10120__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08462_ _03307_ _03321_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07676__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07413_ _02535_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__or2_4
XANTENNA__06884__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08393_ _02635_ _02683_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07344_ top.a1.instruction\[29\] net528 _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06393__X _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06636__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07275_ _02380_ _02399_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout313_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09014_ _03836_ _03852_ _04075_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__or3_1
XANTENNA__10983__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06226_ net1890 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[2\] sky130_fd_sc_hd__and2_1
XFILLER_0_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08389__B1 _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold120 top.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
X_06157_ net903 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XANTENNA__10790__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 top.a1.row2\[10\] vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 top.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 top.DUT.register\[8\]\[16\] vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 top.ramload\[28\] vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 top.DUT.register\[23\]\[22\] vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 top.ramstore\[21\] vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout600 _01669_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_2
Xhold197 top.DUT.register\[10\]\[30\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 _01666_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11187__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout622 _01663_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
X_09916_ net145 net1924 net438 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__mux2_1
Xfanout633 net634 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_4
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout644 _01647_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 _01639_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout666 _01636_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_2
XANTENNA__09880__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout677 _01549_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_4
X_09847_ _04844_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nand2_1
Xfanout688 _01543_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 _01537_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout947_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _04394_ net527 net333 top.a1.dataIn\[17\] _04783_ vssd1 vssd1 vccd1 vccd1
+ _04784_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_161_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _02079_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11740_ _05549_ _05572_ _05605_ _05606_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__o32a_1
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07667__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06875__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _05518_ _05521_ _05509_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13410_ clknet_leaf_43_clk _00974_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10622_ net219 net2100 net392 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07419__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13341_ clknet_leaf_104_clk _00905_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _04711_ net2212 net359 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_94_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13272_ clknet_leaf_13_clk _00836_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10484_ net256 net1838 net365 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__mux2_1
X_12223_ _06037_ net590 _06061_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07052__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _06009_ _06011_ _06016_ _06004_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o31a_1
X_11105_ net2127 net857 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__and2_1
XANTENNA__10205__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ _05944_ _05946_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__nor2_1
X_11036_ net16 net842 net812 net1635 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__o22a_1
XANTENNA__11151__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12987_ clknet_leaf_59_clk _00551_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09789__X _04794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__inv_2
XANTENNA__08855__A1 _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12429__Q top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10875__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ _05695_ net131 _05697_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13608_ clknet_leaf_83_clk net1215 net1013 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10447__Y _04958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06618__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ clknet_leaf_41_clk _01103_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07060_ top.a1.instruction\[2\] _01494_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_70_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07291__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06397__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10115__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ _01973_ _01991_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__nand2b_1
X_09701_ _02198_ _02203_ _04151_ _02192_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__and4b_1
X_06913_ top.DUT.register\[30\]\[21\] net715 net688 top.DUT.register\[1\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
X_07893_ top.DUT.register\[20\]\[17\] net576 net627 top.DUT.register\[9\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09632_ _04643_ _04648_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__nor2_1
X_06844_ top.DUT.register\[8\]\[23\] net568 net552 top.DUT.register\[7\]\[23\] _01957_
+ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a221o_1
XANTENNA__06388__X _01515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07897__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _04596_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__nand2_1
X_06775_ top.DUT.register\[10\]\[25\] net600 net541 top.DUT.register\[22\]\[25\] _01901_
+ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08514_ net320 _03628_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09699__X _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08846__A1 _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07649__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ top.pc\[26\] _04515_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06857__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ _03455_ _03562_ net304 vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout430_A _04920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07327_ top.DUT.register\[4\]\[8\] net767 net674 top.DUT.register\[18\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XANTENNA__11602__B1 top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09271__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07282__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07258_ top.DUT.register\[9\]\[14\] net628 net621 top.DUT.register\[26\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07821__A2 _02947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06209_ net890 _01426_ net34 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__o21a_1
X_07189_ _02300_ _02302_ _02306_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__nor4_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13300__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__A1 _02709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _04920_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_4
Xfanout441 _04965_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_8
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 _01625_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
Xfanout485 _03179_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_4
X_12910_ clknet_leaf_117_clk _00474_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07888__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ net1140 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
X_12841_ clknet_leaf_3_clk _00405_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06560__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12772_ clknet_leaf_40_clk _00336_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_169_Left_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11723_ top.a1.dataIn\[9\] _05560_ _05590_ _05591_ vssd1 vssd1 vccd1 vccd1 _05593_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06848__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11654_ _05500_ _05516_ _05520_ _05489_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ net165 net1726 net387 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09798__C1 _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire820 _01575_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_1
X_11585_ _05441_ _05442_ _05432_ _05434_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_181_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ clknet_leaf_9_clk _00888_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10536_ net1448 net183 net364 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__mux2_1
XANTENNA__07812__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13255_ clknet_leaf_6_clk _00819_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_178_Left_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ net205 net2034 net371 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07025__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ _05846_ _04976_ net845 top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 _01291_
+ sky130_fd_sc_hd__a2bb2o_1
X_13186_ clknet_leaf_42_clk _00750_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07576__A1 top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ net229 net2258 net328 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__mux2_1
XANTENNA__08773__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _05993_ _06002_ _06006_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09009__B _03768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12893__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ _05890_ _05907_ _05896_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_205_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11019_ net29 net832 net830 net2342 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__a22o_1
XANTENNA__07879__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06551__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06560_ top.DUT.register\[12\]\[30\] net608 net596 top.DUT.register\[27\]\[30\] _01675_
+ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06491_ top.a1.instruction\[2\] _01494_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__and2_4
XFILLER_0_75_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06303__A2 _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08230_ _03217_ _03241_ net279 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08161_ _03284_ _03286_ net282 vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07112_ top.DUT.register\[3\]\[12\] net690 net669 top.DUT.register\[5\]\[12\] _02238_
+ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a221o_1
X_08092_ _03211_ _03218_ net302 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07264__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07803__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload40 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload40/X sky130_fd_sc_hd__clkbuf_8
X_07043_ top.DUT.register\[27\]\[10\] net775 net685 top.DUT.register\[1\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
Xclkload51 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload62 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__clkinv_8
Xclkload73 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload73/X sky130_fd_sc_hd__clkbuf_8
Xclkload84 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload95 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_8
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08104__A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ _03717_ _03739_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1018_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _03068_ _03069_ _03070_ _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_145_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_A _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06790__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ top.DUT.register\[21\]\[17\] net692 net671 top.DUT.register\[16\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_1
X_09615_ top.pad.keyCode\[4\] top.pad.keyCode\[6\] top.pad.keyCode\[7\] top.pad.keyCode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__or4b_2
X_06827_ top.DUT.register\[22\]\[23\] net751 net678 top.DUT.register\[13\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout645_A _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ _04575_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__and2_1
X_06758_ _01875_ _01880_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__nor3_1
XFILLER_0_210_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ top.pc\[24\] _04483_ top.pc\[25\] vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_191_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06689_ net807 _01815_ _01624_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09492__B2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08428_ _02587_ _03516_ _03525_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
X_08359_ _02634_ _03177_ net483 _02635_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09809__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07255__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11370_ _05223_ _05224_ _05211_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10321_ net1724 net214 net399 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07007__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ clknet_leaf_0_clk _00604_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10252_ net1478 net211 net457 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__mux2_1
X_10183_ net228 net1639 net412 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
XANTENNA__10562__A0 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08949__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input39_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 net262 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
Xfanout271 _03238_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
Xfanout282 _02856_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
Xfanout293 _02811_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12434__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06469__A top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13873_ net1160 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_202_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12824_ clknet_leaf_13_clk _00388_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13541__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ clknet_leaf_1_clk _00319_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09483__A1 _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11706_ _05534_ _05575_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07494__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12686_ clknet_leaf_118_clk _00250_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11637_ _05473_ _05501_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07246__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06491__X _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ _05437_ _05404_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_188_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ clknet_leaf_57_clk _00871_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold708 top.DUT.register\[2\]\[30\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold719 top.DUT.register\[31\]\[21\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ net1802 net248 net361 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__mux2_1
X_11499_ _05322_ _05368_ _05365_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13238_ clknet_leaf_120_clk _00802_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12442__Q top.a1.dataIn\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10553__A0 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ clknet_leaf_12_clk _00733_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07763__A _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06772__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07730_ top.DUT.register\[27\]\[1\] net777 net745 top.DUT.register\[31\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07661_ net529 _02424_ _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__a21bo_4
XTAP_TAPCELL_ROW_0_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ net512 _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and2b_1
X_06612_ top.DUT.register\[24\]\[28\] net738 net722 top.DUT.register\[14\]\[28\] _01738_
+ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ top.DUT.register\[27\]\[3\] net775 net689 top.DUT.register\[3\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
X_09331_ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__inv_2
X_06543_ _01590_ _01630_ _01643_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__and3_4
XANTENNA__09474__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06385__Y _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09262_ net894 _04304_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__and2_1
XANTENNA__11281__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06474_ top.a1.instruction\[7\] top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 _01601_
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08213_ _03161_ _03173_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09193_ _04233_ _04237_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout226_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08144_ _03268_ _03269_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__nand2_1
XANTENNA__07237__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11033__B2 top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08075_ net296 _03127_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09787__A1_N net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07026_ top.DUT.register\[6\]\[11\] net559 net629 top.DUT.register\[9\]\[11\] _02152_
+ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout595_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 _01369_ vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10370__Y _04945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold24 _01175_ vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net1321 net865 _01815_ net593 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__a22o_1
Xhold35 top.ramstore\[6\] vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A _01510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 top.ramstore\[11\] vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06763__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 net92 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ top.DUT.register\[19\]\[16\] net632 net786 top.DUT.register\[3\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__a22o_1
Xhold68 _01187_ vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 top.ramstore\[18\] vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _02977_ _02979_ _02981_ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ net2297 net149 net345 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08981__A1_N _03146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ net910 top.pc\[27\] _04565_ net897 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_158_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06736__B _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12540_ clknet_leaf_93_clk _00104_ net999 vssd1 vssd1 vccd1 vccd1 top.pc\[23\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07476__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__X _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ clknet_leaf_97_clk top.ru.next_FetchedInstr\[23\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[23\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_193_Right_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11422_ _05289_ _05290_ _05261_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07228__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09768__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08976__B1 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__B2 _02143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ _05217_ _05219_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_104_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06471__B top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10304_ net1694 net263 net398 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11284_ top.a1.row1\[60\] _05112_ _01444_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13023_ clknet_leaf_113_clk _00587_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09782__B _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10235_ net1751 net264 net456 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__mux2_1
Xfanout1000 net1020 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07583__A _02709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07400__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1022 net1029 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
X_10166_ net464 _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__nand2_1
Xfanout1033 net1038 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06754__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 net1051 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
Xfanout1055 net1060 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_2
Xfanout1077 net1079 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10213__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06199__A top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10097_ _01601_ _04676_ _04921_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__nor3_1
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1099 net1102 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload4_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13856_ net1121 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XANTENNA__06486__X _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12807_ clknet_leaf_26_clk _00371_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13787_ clknet_leaf_67_clk _01330_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10999_ top.a1.dataIn\[8\] net848 net843 _05014_ vssd1 vssd1 vccd1 vccd1 _05015_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11263__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ clknet_leaf_43_clk _00302_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07467__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13403__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__B2 top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10883__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12669_ clknet_leaf_105_clk _00233_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07219__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06190_ _01411_ _01418_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__nand2_2
XANTENNA__12212__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08967__B1 _03031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold505 top.DUT.register\[12\]\[31\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 top.DUT.register\[25\]\[6\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__A2 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06381__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 top.DUT.register\[11\]\[0\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold538 top.DUT.register\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 top.DUT.register\[7\]\[5\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08900_ _01735_ _03978_ _01734_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o21bai_1
X_09880_ net833 _04555_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08831_ net268 _03373_ _03878_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_5_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06745__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ _02037_ _03850_ _02035_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a21oi_1
X_07713_ top.DUT.register\[17\]\[1\] net645 net621 top.DUT.register\[26\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a22o_1
X_08693_ _03764_ _03800_ net280 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout176_A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ _02763_ _02765_ _02767_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06396__X _01523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07575_ top.DUT.register\[19\]\[3\] net631 net779 top.DUT.register\[15\]\[3\] _02692_
+ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a221o_1
X_09314_ _02331_ _02338_ _04362_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__or3_2
XFILLER_0_180_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06526_ _01628_ _01631_ _01637_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__and3_4
XFILLER_0_158_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09245_ _04296_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__nor2_1
XANTENNA__10793__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06457_ net902 _01388_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout608_A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12203__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ _02562_ _02566_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nand2_1
X_06388_ _01497_ _01498_ net790 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__and3_4
XFILLER_0_16_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ net268 _03236_ net272 _03253_ _03222_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a221o_1
X_08058_ net277 _03168_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_186_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06984__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A2 _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ _02132_ _02133_ _02135_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__or3_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
X_10020_ net178 top.DUT.register\[4\]\[23\] net425 vssd1 vssd1 vccd1 vccd1 _00241_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09922__A2 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10033__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _05817_ _05826_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13710_ clknet_leaf_72_clk _01258_ net1096 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_98_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10922_ net203 net2174 net444 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XANTENNA__07697__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07161__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13641_ clknet_leaf_83_clk _01200_ net1011 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10853_ net2135 net229 net350 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13641__Q net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06466__B top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ clknet_leaf_84_clk _01131_ net1017 vssd1 vssd1 vccd1 vccd1 top.a1.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10784_ net1848 net202 net447 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12523_ clknet_leaf_78_clk _00087_ net1003 vssd1 vssd1 vccd1 vccd1 top.pc\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ clknet_leaf_100_clk top.ru.next_FetchedInstr\[6\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06482__A top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ _05244_ _05256_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__nand2b_1
X_12385_ clknet_leaf_88_clk _00021_ net1006 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10208__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__A1 _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11336_ top.a1.dataIn\[20\] _05189_ _05193_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__and3_1
XANTENNA__07621__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06975__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ top.a1.row1\[106\] _05116_ _05119_ top.a1.row1\[18\] _05144_ vssd1 vssd1
+ vccd1 vccd1 _05145_ sky130_fd_sc_hd__a221o_1
X_13006_ clknet_leaf_111_clk _00570_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10218_ net215 net2299 net405 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_105_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11198_ net1237 _05079_ _05086_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__a21o_1
XANTENNA__06727__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09017__B _03606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ net229 net1313 net414 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10878__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__B2 top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__B _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07688__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07105__X _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09033__A _03715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ net72 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11713__D top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ top.DUT.register\[28\]\[8\] net651 net599 top.DUT.register\[10\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_114_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06311_ _01451_ _01332_ _01452_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__nand3_1
X_07291_ top.DUT.register\[9\]\[9\] net711 net697 top.DUT.register\[23\]\[9\] _02416_
+ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ _03798_ _03914_ _03926_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__and4_1
XFILLER_0_170_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06242_ net1386 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[18\] sky130_fd_sc_hd__and2_1
XANTENNA__07860__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06173_ top.pad.button_control.r_counter\[8\] vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XANTENNA__10118__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12537__RESET_B net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold302 top.DUT.register\[23\]\[3\] vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 top.DUT.register\[3\]\[29\] vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 top.DUT.register\[22\]\[9\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09907__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold335 top.DUT.register\[11\]\[29\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 top.DUT.register\[7\]\[3\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 top.DUT.register\[29\]\[30\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 top.DUT.register\[13\]\[26\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net253 net1793 net435 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold379 top.DUT.register\[30\]\[8\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 _01585_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07778__A_N _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__B1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout815 net818 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_2
XFILLER_0_111_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout826 net827 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_2
XANTENNA__09208__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ top.pc\[26\] _04543_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__nand2_1
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_2
XANTENNA__08112__A _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_A _02811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_181_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _03898_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__nand2_1
Xhold1002 top.DUT.register\[10\]\[12\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 top.DUT.register\[13\]\[30\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 top.DUT.register\[27\]\[6\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09794_ _04787_ _04790_ _04796_ _01586_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a31o_1
Xhold1035 top.DUT.register\[29\]\[14\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 top.DUT.register\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 top.DUT.register\[7\]\[8\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ _03817_ _03849_ _02077_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout460_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__A1 _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 top.DUT.register\[21\]\[25\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 top.DUT.register\[15\]\[20\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout558_A _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ net315 _03374_ _03543_ net478 vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_200_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07015__X _02142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08340__B2 _03462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ _02746_ _02748_ _02750_ _02753_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_132_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout725_A _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07558_ _02683_ _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__nand2_2
XFILLER_0_76_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06509_ _01591_ net789 _01634_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08643__A2 _03741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__A1 _03882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ top.DUT.register\[14\]\[5\] net611 net595 top.DUT.register\[27\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ _04280_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__or2_1
XANTENNA__07851__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09159_ _02642_ _02682_ _04206_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_133_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10028__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ _06035_ _06036_ _06034_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_141_Left_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06957__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ net52 net859 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__and2_1
Xhold880 top.DUT.register\[20\]\[4\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold891 top.DUT.register\[17\]\[8\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_166_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ net98 net856 net825 net1175 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08022__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ net245 net1229 net427 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10698__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06590__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ _05822_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_Left_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07134__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ net260 net1649 net441 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
X_11885_ _05702_ _05738_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13624_ clknet_leaf_75_clk net1257 net1088 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10836_ net464 _04940_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_15_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13555_ clknet_leaf_68_clk _01119_ net1104 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ net157 net1784 net376 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ clknet_leaf_45_clk _00073_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramstore\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13486_ clknet_leaf_115_clk _01050_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10698_ net176 net1745 net377 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12437_ clknet_leaf_94_clk top.ru.next_FetchedData\[21\] net995 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[21\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__12194__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09595__B1 _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ top.pad.button_control.r_counter\[15\] _06148_ vssd1 vssd1 vccd1 vccd1 _06151_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ _05186_ _05187_ _05188_ _05184_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12299_ top.lcd.cnt_500hz\[7\] _06106_ _06098_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_130_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09028__A _03619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13836__RESET_B net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06860_ top.DUT.register\[9\]\[23\] net708 net671 top.DUT.register\[16\]\[23\] _01986_
+ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a221o_1
XANTENNA__07373__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ top.DUT.register\[12\]\[24\] net582 net672 top.DUT.register\[16\]\[24\] _01910_
+ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a221o_1
XANTENNA__06581__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08530_ _03643_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10401__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08322__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07125__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08461_ _03577_ _03578_ net317 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07412_ _02525_ _02536_ _02537_ _02538_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__or4_1
X_08392_ net519 _03503_ _03512_ net479 _03510_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_34_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07343_ _02185_ _02424_ _02207_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07833__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ _02400_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__inv_2
X_09013_ _03799_ _03932_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06225_ net2102 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[1\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout306_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__A1 _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 _01186_ vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08389__B2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 net94 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ net906 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold132 top.DUT.register\[20\]\[9\] vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 top.ramaddr\[9\] vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 top.DUT.register\[24\]\[18\] vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 top.ramload\[27\] vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 top.ramstore\[17\] vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_8
Xhold187 top.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _01666_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_2
Xhold198 top.ramaddr\[31\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ net336 _04901_ _04907_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__and3_2
Xfanout623 _01662_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_8
Xfanout634 _01656_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XANTENNA_fanout675_A _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _01647_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout656 _01639_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
X_09846_ top.pc\[24\] _04508_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__or2_1
Xfanout667 _01554_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08010__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net680 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_8
Xfanout689 net691 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ net834 _04387_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nor2_1
X_06989_ top.DUT.register\[8\]\[20\] net570 net553 top.DUT.register\[7\]\[20\] _02105_
+ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06572__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _02119_ _03817_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__and2b_1
XANTENNA__10311__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__A2 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ net522 _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11670_ _05533_ _05538_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10621_ net225 net1661 net390 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09895__X _04890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ clknet_leaf_77_clk _00904_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10552_ net246 net1770 net357 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__Q top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13271_ clknet_leaf_106_clk _00835_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10483_ net262 net1826 net365 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12222_ net1192 net590 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _06011_ _06016_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ net916 net1306 net853 _05038_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a31o_1
XANTENNA__11097__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ _05949_ _05952_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__or3_1
XANTENNA__07862__Y _02989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ net15 net831 net830 top.ramload\[21\] vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__a22o_1
XANTENNA__08001__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__B2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10221__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ clknet_leaf_15_clk _00550_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11937_ _05803_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__nor2_1
XANTENNA__08855__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11868_ _05695_ _05697_ net131 vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and3_1
XFILLER_0_200_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ clknet_leaf_92_clk _01166_ net1000 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_2
X_10819_ net1379 net181 net353 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__mux2_1
X_11799_ _05613_ _05665_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_119_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07815__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13538_ clknet_leaf_41_clk _01102_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10891__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13469_ clknet_leaf_103_clk _01033_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08791__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__B2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ net512 _02118_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__and2b_1
X_09700_ net241 net1757 net438 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06912_ top.DUT.register\[16\]\[21\] _01514_ net699 top.DUT.register\[23\]\[21\]
+ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a221o_1
X_07892_ top.DUT.register\[7\]\[17\] net552 net603 top.DUT.register\[18\]\[17\] _03018_
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__a221o_1
XANTENNA__07346__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _04644_ _04647_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11142__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06843_ top.DUT.register\[11\]\[23\] net639 net548 top.DUT.register\[24\]\[23\] _01958_
+ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a221o_1
XANTENNA__06554__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ top.pc\[29\] _04578_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__or2_1
X_06774_ top.DUT.register\[17\]\[25\] net644 net624 top.DUT.register\[25\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08513_ net274 _03398_ _03406_ net270 vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__o22a_1
X_09493_ _04524_ _04531_ top.pc\[25\] _04044_ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_188_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08444_ _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08536__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ _03293_ _03409_ _03495_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout423_A _04925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07326_ top.DUT.register\[1\]\[8\] net685 net678 top.DUT.register\[13\]\[8\] _02452_
+ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07806__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09875__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07257_ top.DUT.register\[1\]\[14\] net657 net641 top.DUT.register\[11\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06208_ top.ru.state\[2\] top.busy_o vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__and2_1
X_07188_ _02308_ _02310_ _02312_ _02314_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07395__B net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10306__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 _04927_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
XANTENNA__06793__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__Y _03882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 net432 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
Xfanout442 _04965_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
Xfanout453 _04946_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_8
Xfanout464 _04677_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_12
XANTENNA__07337__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 net477 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 _03179_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
X_09829_ net802 _04826_ _04827_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a31o_1
XANTENNA__06545__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ clknet_leaf_32_clk _00404_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10041__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ clknet_leaf_22_clk _00335_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11722_ _05590_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08446__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09131__A _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11653_ _05517_ _05518_ _05521_ _05490_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__o31a_1
XFILLER_0_153_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09798__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ net169 net2228 net388 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11584_ _05441_ _05442_ _05434_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ clknet_leaf_29_clk _00887_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10535_ net1605 net189 net364 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08470__B1 _03584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ clknet_leaf_25_clk _00818_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10466_ net212 net1952 net372 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12205_ top.a1.row2\[32\] net845 net813 net127 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__a22o_1
XANTENNA__10216__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ clknet_leaf_27_clk _00749_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10397_ net180 net1603 net328 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__mux2_1
XANTENNA__07576__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12136_ _05981_ _05985_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09009__C _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06784__B1 _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ _05933_ _05936_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__nand2_1
XANTENNA__07328__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output52_A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net28 net841 net811 net1553 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__o22a_1
XANTENNA__09722__B1 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10886__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ clknet_leaf_11_clk _00533_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06490_ net821 _01615_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07500__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09238__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08160_ _01840_ net292 _03285_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_172_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ top.DUT.register\[25\]\[12\] net774 net765 top.DUT.register\[6\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08091_ _03214_ _03217_ net276 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload30 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__bufinv_16
Xclkload41 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload41/X sky130_fd_sc_hd__clkbuf_4
X_07042_ top.DUT.register\[20\]\[10\] net748 _01535_ top.DUT.register\[3\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload52 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__clkinv_4
Xclkload63 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__inv_6
Xclkload74 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload85 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload85/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10126__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload96 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_16
XANTENNA__10020__A0 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _03666_ _03673_ _03711_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_54_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06775__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__A top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07944_ top.DUT.register\[20\]\[16\] net577 net608 top.DUT.register\[12\]\[16\] _03056_
+ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_145_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09216__A _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__A _02143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _02997_ _02999_ _03000_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__or4_4
XFILLER_0_207_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout373_A _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ top.pad.keyCode\[1\] top.pad.keyCode\[0\] top.pad.keyCode\[2\] top.pad.keyCode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__or4b_4
X_06826_ _01950_ _01951_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_178_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _04579_ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06757_ _01881_ _01882_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__or3_1
XANTENNA__10796__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout540_A _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12733__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ top.pc\[24\] top.pc\[25\] _04483_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ top.DUT.register\[20\]\[27\] net576 _01812_ _01813_ _01814_ vssd1 vssd1 vccd1
+ vccd1 _01815_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08427_ net519 _03546_ _03540_ _03539_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout805_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08358_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload2 clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_22_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07309_ top.DUT.register\[20\]\[9\] net577 _02433_ _02435_ vssd1 vssd1 vccd1 vccd1
+ _02436_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08289_ net312 _02731_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_210_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ top.DUT.register\[13\]\[17\] net215 net397 vssd1 vssd1 vccd1 vccd1 _00523_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ net1456 net217 net454 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10036__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net179 net2220 net409 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
Xfanout250 _05407_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_1
XANTENNA__11106__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 _03237_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xfanout283 _02712_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XANTENNA__13644__Q net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__D_N _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13872_ net1159 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_202_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12823_ clknet_leaf_17_clk _00387_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10078__A0 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ clknet_leaf_53_clk _00318_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11705_ _05533_ _05559_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12685_ clknet_leaf_22_clk _00249_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11290__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11636_ _05478_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11567_ _05399_ net250 vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07797__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ net1446 net254 net363 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ clknet_leaf_17_clk _00870_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 top.DUT.register\[13\]\[3\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _05339_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or2_2
XANTENNA__08205__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13237_ clknet_leaf_6_clk _00801_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10449_ net265 net2093 net371 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__09943__A0 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ clknet_leaf_122_clk _00732_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _05987_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__nor2_1
X_13099_ clknet_leaf_23_clk _00663_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11285__B _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07660_ _02209_ _02785_ _02207_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XANTENNA__07182__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13366__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ top.DUT.register\[26\]\[28\] net762 net698 top.DUT.register\[23\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07591_ top.DUT.register\[26\]\[3\] net759 net692 top.DUT.register\[21\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _01615_ _02610_ _02638_ net821 _01622_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_149_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06542_ _01631_ _01637_ _01643_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__and3_4
XFILLER_0_48_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07485__A1 top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _04298_ _04300_ _04297_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a21o_1
X_06473_ top.a1.instruction\[3\] top.a1.instruction\[6\] top.a1.instruction\[15\]
+ top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_173_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08682__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08212_ _03161_ _03173_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__and2_2
XFILLER_0_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09192_ _02516_ _02521_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ net514 net292 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout219_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _01560_ net296 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08115__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07025_ top.DUT.register\[16\]\[11\] net638 net598 top.DUT.register\[27\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08737__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06212__A2 top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ net1241 net869 _01858_ net594 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a22o_1
Xhold25 top.ramstore\[10\] vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _01173_ vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _01178_ vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 _01194_ vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _03045_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__nor2_8
XFILLER_0_194_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold69 top.DUT.register\[4\]\[6\] vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_A _01515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07858_ top.DUT.register\[13\]\[18\] net650 net629 top.DUT.register\[9\]\[18\] _02984_
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a221o_1
XANTENNA__07173__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07712__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06809_ top.DUT.register\[20\]\[24\] net578 net566 top.DUT.register\[4\]\[24\] _01935_
+ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ top.DUT.register\[23\]\[19\] net698 net683 top.DUT.register\[7\]\[19\] _02915_
+ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a221o_1
XFILLER_0_210_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06920__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11257__C1 _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ net132 _04554_ _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08963__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ net136 _04485_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_80_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12470_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[22\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[22\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11421_ _05289_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08978__A2_N net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08976__B2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ top.a1.dataIn\[29\] top.a1.dataIn\[30\] _05194_ vssd1 vssd1 vccd1 vccd1 _05222_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06987__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06471__C top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net1557 net150 net397 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11283_ net1225 net824 _05159_ net1091 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__o211a_1
X_13022_ clknet_leaf_14_clk _00586_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10234_ net1687 net150 net454 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__mux2_1
XANTENNA__07864__A _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06739__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__B1 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
X_10165_ _04679_ _04929_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1023 net1029 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_210_Right_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1034 net1038 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13389__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1045 net1050 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 net1060 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__clkbuf_4
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_2
X_10096_ net140 net2186 net419 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1089 net1092 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13855_ net1120 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XANTENNA__06911__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12806_ clknet_leaf_24_clk _00370_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13786_ clknet_leaf_64_clk _01329_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10998_ top.a1.data\[4\] top.a1.dataInTemp\[8\] net797 vssd1 vssd1 vccd1 vccd1 _05014_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09797__Y _04801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ clknet_leaf_26_clk _00301_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08664__B1 _03763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A2 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12668_ clknet_leaf_17_clk _00232_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12212__A1 top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _05446_ _05485_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12599_ clknet_leaf_106_clk _00163_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08967__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold506 top.DUT.register\[31\]\[17\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06978__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire492 _03126_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12453__Q top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold517 top.DUT.register\[18\]\[16\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold528 top.DUT.register\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 top.DUT.register\[3\]\[26\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ net316 _03605_ _03788_ _03237_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_51_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10404__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08761_ net1279 net837 net816 _03865_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a22o_1
XANTENNA__12756__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ top.DUT.register\[4\]\[1\] net566 net563 top.DUT.register\[23\]\[1\] _02838_
+ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a221o_1
X_08692_ _03272_ _03276_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__nand2_1
X_13860__1151 vssd1 vssd1 vccd1 vccd1 net1151 _13860__1151/LO sky130_fd_sc_hd__conb_1
XANTENNA__07155__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07643_ top.DUT.register\[31\]\[2\] net743 net735 top.DUT.register\[24\]\[2\] _02761_
+ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout169_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07574_ top.DUT.register\[4\]\[3\] net564 net615 top.DUT.register\[30\]\[3\] _02700_
+ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09313_ _01615_ _02638_ _02688_ net823 _01622_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__o221a_2
XFILLER_0_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06525_ _01632_ _01651_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_196_Left_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout336_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09244_ _02212_ top.pc\[11\] vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__and2b_1
X_06456_ _01478_ _01479_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07949__A _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09175_ _02562_ _02566_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_153_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06387_ _01496_ net793 _01505_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__and3_4
XANTENNA__06681__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12203__B2 top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _03245_ _03252_ net302 vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__mux2_1
XANTENNA__08958__B2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08057_ _03172_ _03182_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_186_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07008_ top.DUT.register\[14\]\[11\] net722 net703 top.DUT.register\[29\]\[11\] _02134_
+ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__10381__Y _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_168_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10314__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09922__A3 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ net501 net591 net1190 net867 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _05831_ _05835_ _05837_ _05839_ _05808_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_169_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10921_ net211 net1621 net443 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
X_10852_ net1408 net182 net350 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
X_13640_ clknet_leaf_88_clk _01199_ net1006 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12538__Q top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06466__C top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ clknet_leaf_84_clk _01130_ net1015 vssd1 vssd1 vccd1 vccd1 top.a1.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10783_ net1427 net209 net447 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12522_ clknet_leaf_78_clk _00086_ net1004 vssd1 vssd1 vccd1 vccd1 top.pc\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12453_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[5\] net997 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[5\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__06672__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ _05199_ _05227_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12384_ clknet_leaf_82_clk _00020_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11335_ top.a1.dataIn\[21\] _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06424__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11266_ top.a1.row2\[10\] _05117_ _05118_ top.a1.row2\[18\] vssd1 vssd1 vccd1 vccd1
+ _05144_ sky130_fd_sc_hd__a22o_1
XANTENNA__09374__A1 top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ net228 net1645 net406 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__mux2_1
X_13005_ clknet_leaf_33_clk _00569_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10224__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ net850 _05072_ net531 vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__and3_1
XANTENNA__07385__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net180 net1733 net413 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
XANTENNA__09126__A1 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ net196 net2104 net419 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__mux2_1
XANTENNA__07137__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ net72 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10894__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ clknet_leaf_65_clk _01312_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_42_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06310_ _01332_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07290_ top.DUT.register\[31\]\[9\] net743 net692 top.DUT.register\[21\]\[9\] _02414_
+ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a221o_1
XANTENNA__08217__X _03343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06241_ net1333 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[17\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12197__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06172_ net1172 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__A1_N net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold303 top.a1.row1\[120\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08808__A2_N net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold314 top.DUT.register\[21\]\[15\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 top.DUT.register\[7\]\[18\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06415__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 top.DUT.register\[7\]\[24\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 top.DUT.register\[28\]\[13\] vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold358 top.DUT.register\[19\]\[28\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 top.DUT.register\[23\]\[21\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net256 net1959 net433 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_3__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout805 net807 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout816 net817 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_7__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_1
X_09862_ top.pc\[25\] _04518_ _04853_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09208__B _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08887__X _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout838 net840 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07376__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout849 _04634_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07915__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1003 top.DUT.register\[30\]\[10\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net474 _03902_ _03914_ net471 _03912_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_181_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09793_ _04787_ _04790_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a21oi_1
Xhold1014 top.DUT.register\[31\]\[19\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 top.DUT.register\[28\]\[18\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09117__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1036 top.DUT.register\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 top.DUT.register\[10\]\[14\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07951__B _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1058 top.DUT.register\[26\]\[19\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _02078_ _02119_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__nor2_1
XANTENNA__09668__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 top.DUT.register\[18\]\[1\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _02993_ _03083_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ top.DUT.register\[7\]\[2\] net552 net615 top.DUT.register\[30\]\[2\] _02752_
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a221o_1
XFILLER_0_191_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ net319 _02682_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout620_A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06508_ _01628_ net789 _01634_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__and3_4
XFILLER_0_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07488_ top.DUT.register\[23\]\[5\] net560 net548 top.DUT.register\[24\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06439_ top.a1.instruction\[0\] top.a1.instruction\[1\] top.a1.instruction\[2\] vssd1
+ vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__and3_1
XANTENNA__06654__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09227_ top.pc\[9\] _04254_ top.pc\[10\] vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10309__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09158_ _04213_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08109_ net306 _03233_ _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__o21ai_1
X_09089_ _02193_ _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ net915 net1332 net853 _05046_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08303__A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 top.ru.state\[6\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 top.DUT.register\[27\]\[30\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 top.DUT.register\[5\]\[17\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net1254 net856 net825 top.ramstore\[2\] vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a22o_1
XANTENNA__10044__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10002_ net247 net1725 net425 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07119__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _05786_ _05789_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nand2_4
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10904_ net264 net1438 net443 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ _05745_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_196_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13623_ clknet_leaf_83_clk net1178 net1014 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06893__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ net2348 net142 net355 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_15_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13554_ clknet_leaf_69_clk _01118_ net1104 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ net162 net1655 net373 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ clknet_leaf_45_clk _00072_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramstore\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06645__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10219__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697_ net184 net2221 net380 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ clknet_leaf_23_clk _01049_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12436_ clknet_leaf_94_clk top.ru.next_FetchedData\[20\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12367_ top.pad.button_control.r_counter\[15\] _06148_ vssd1 vssd1 vccd1 vccd1 _06150_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11318_ top.a1.dataIn\[23\] top.a1.dataIn\[21\] top.a1.dataIn\[20\] top.a1.dataIn\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__or4bb_1
X_12298_ _06106_ _06098_ _06105_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_130_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11249_ net1219 net824 _05128_ net1093 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__o211a_1
XANTENNA_max_cap516_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10889__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07771__B _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ top.DUT.register\[9\]\[24\] net709 net687 top.DUT.register\[1\]\[24\] _01916_
+ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_11__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__08858__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ net311 _03349_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07411_ top.DUT.register\[21\]\[7\] net573 net599 top.DUT.register\[10\]\[7\] _02524_
+ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08391_ net319 _03511_ _03502_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11209__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07342_ _02458_ _02460_ _02468_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__nor3_1
XFILLER_0_9_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08094__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ _02380_ _02399_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__and2_1
XANTENNA__10129__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _03475_ _03503_ _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__nand4_1
X_06224_ net1340 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[0\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08389__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 net81 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06155_ top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout201_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold111 top.ramaddr\[13\] vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _01196_ vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold133 top.a1.row1\[104\] vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 top.ramaddr\[5\] vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold155 top.ramaddr\[4\] vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08123__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 top.a1.row2\[1\] vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 top.DUT.register\[3\]\[30\] vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 top.pad.button_control.r_counter\[12\] vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold199 top.ramload\[3\] vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _04903_ _04904_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout602 _01669_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_8
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_4
XANTENNA__07349__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 _01662_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1110_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 _01652_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_4
Xfanout646 _01647_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ top.pc\[24\] _04508_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nand2_1
Xfanout657 _01639_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10799__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _01554_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_2
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout668_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ net802 _04779_ _04781_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__and3_1
X_06988_ _02107_ _02109_ _02111_ _02114_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__or4_1
X_08727_ net1312 net837 net816 _03833_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__a22o_1
XANTENNA__06297__B _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12545__SET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ net274 _03766_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07521__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__D net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07609_ net901 net524 _02735_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_194_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06875__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ _03603_ _03701_ net304 vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09401__B net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ net233 net1484 net390 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ net254 net2040 net359 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__mux2_1
XANTENNA__10039__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09026__B1 _03741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ clknet_leaf_121_clk _00834_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10482_ net265 net2229 net367 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__mux2_1
XANTENNA__12499__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11659__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ net1179 _06045_ net589 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07588__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _05990_ _06013_ _06018_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a31oi_1
XANTENNA__07052__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11103_ net42 net860 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12083_ _05928_ _05950_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__xnor2_4
XANTENNA__11136__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ net14 net841 net811 net2156 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__o22a_1
X_13854__1119 vssd1 vssd1 vccd1 vccd1 _13854__1119/HI net1119 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_188_Right_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08552__A2 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ clknet_leaf_34_clk _00549_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11936_ _05776_ _05786_ _05790_ _05781_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_59_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11867_ _05695_ net131 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13606_ clknet_leaf_98_clk _01165_ net981 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07768__A_N net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10818_ net1319 net197 net355 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__mux2_1
XANTENNA__11292__C_N top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ _05606_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_119_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06618__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ clknet_leaf_27_clk _01101_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10749_ net225 top.DUT.register\[26\]\[10\] net374 vssd1 vssd1 vccd1 vccd1 _00932_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07291__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06951__A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13468_ clknet_leaf_53_clk _01032_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12419_ clknet_leaf_96_clk top.ru.next_FetchedData\[3\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07579__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ clknet_leaf_17_clk _00963_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__Q top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08791__A2 _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ _02076_ _02056_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_4_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_56_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06911_ top.DUT.register\[25\]\[21\] net773 net729 top.DUT.register\[10\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a22o_1
X_07891_ top.DUT.register\[29\]\[17\] net663 net607 top.DUT.register\[12\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09630_ _04652_ _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__or2_1
X_06842_ _01960_ _01962_ _01964_ _01968_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__or4_1
XANTENNA__09740__B2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10412__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09561_ top.pc\[29\] _04578_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__nand2_1
X_06773_ top.DUT.register\[29\]\[25\] net664 net561 top.DUT.register\[23\]\[25\] _01899_
+ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a221o_1
X_08512_ net284 _03430_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06306__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09492_ net136 _04517_ _04530_ net132 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__o22a_1
XFILLER_0_188_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08443_ _03504_ _03561_ net277 vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__mux2_1
XANTENNA__06857__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout151_A _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout249_A _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08374_ net302 _03371_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_176_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09256__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07325_ top.DUT.register\[31\]\[8\] net743 net716 top.DUT.register\[2\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11063__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1060_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout416_A _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07256_ top.DUT.register\[2\]\[14\] net662 net637 top.DUT.register\[16\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
XANTENNA__07282__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06207_ net874 top.ru.next_dready net34 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__or3b_1
X_07187_ top.DUT.register\[4\]\[13\] net565 net626 top.DUT.register\[25\]\[13\] _02313_
+ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a221o_1
XANTENNA__12521__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout785_A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout410 net412 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_6
XANTENNA__08519__C1 _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 _04925_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_6
Xfanout432 _04920_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_8
Xfanout454 _04936_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _04677_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_4
X_09828_ net834 _04470_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__o21bai_1
Xfanout487 net489 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10322__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ net534 _04152_ _04719_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ clknet_leaf_42_clk _00334_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11721_ top.a1.dataIn\[10\] _05528_ _05559_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06848__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09131__B _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11652_ _05517_ _05518_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13873__1160 vssd1 vssd1 vccd1 vccd1 net1160 _13873__1160/LO sky130_fd_sc_hd__conb_1
X_10603_ net172 net1936 net388 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11583_ _05441_ _05442_ _05424_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13322_ clknet_leaf_38_clk _00886_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10534_ net1454 net191 net364 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08470__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13253_ clknet_leaf_120_clk _00817_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ net216 top.DUT.register\[17\]\[17\] net369 vssd1 vssd1 vccd1 vccd1 _00651_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12204_ _05901_ _04976_ net847 top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 _01289_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07025__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13184_ clknet_leaf_46_clk _00748_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10396_ net195 top.DUT.register\[15\]\[14\] net330 vssd1 vssd1 vccd1 vccd1 _00584_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12135_ _05993_ _06002_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07981__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _05896_ _05932_ _05909_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13468__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ net27 net831 net830 net1359 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__a22o_1
XANTENNA__10232__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07733__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12968_ clknet_leaf_33_clk _00532_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06839__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _05776_ _05783_ _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_169_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12899_ clknet_leaf_22_clk _00463_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09789__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ top.DUT.register\[8\]\[12\] net740 net736 top.DUT.register\[24\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
X_08090_ _03215_ _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__nand2_1
XANTENNA__07264__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload20 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_113_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07041_ top.DUT.register\[24\]\[10\] net735 net716 top.DUT.register\[2\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a22o_1
Xclkload31 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_8
Xclkload42 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload42/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10407__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload53 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload64 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_6
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload75 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_51_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload86 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_140_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload97 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_54_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08992_ _03550_ _03634_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__and3_1
X_07943_ top.DUT.register\[8\]\[16\] net571 net541 top.DUT.register\[22\]\[16\] _03058_
+ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_145_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout199_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09216__B _02427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ top.DUT.register\[27\]\[17\] net775 net689 top.DUT.register\[3\]\[17\] _02995_
+ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a221o_1
XANTENNA__07724__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09931__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ _01604_ _04633_ _04640_ top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1 _00115_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06825_ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout366_A _04959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09544_ _01755_ _04577_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__and2_1
XANTENNA__09477__B1 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06756_ top.DUT.register\[27\]\[25\] net776 net683 top.DUT.register\[7\]\[25\] _01877_
+ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09232__A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__B1 _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13750__Q top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ _04178_ _04507_ _04514_ _04044_ top.pc\[24\] vssd1 vssd1 vccd1 vccd1 _00105_
+ sky130_fd_sc_hd__o32a_1
X_06687_ top.DUT.register\[21\]\[27\] net573 net564 top.DUT.register\[4\]\[27\] _01798_
+ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_191_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ _03532_ _03544_ _03530_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_82_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08357_ net273 _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13853__1118 vssd1 vssd1 vccd1 vccd1 _13853__1118/HI net1118 sky130_fd_sc_hd__conb_1
XANTENNA_fanout700_A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_22_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07308_ top.DUT.register\[28\]\[9\] net652 net616 top.DUT.register\[30\]\[9\] _02434_
+ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07255__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ net314 _03411_ _03402_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08135__X _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10317__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ top.DUT.register\[8\]\[14\] net741 net714 top.DUT.register\[30\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a22o_1
X_10250_ net1390 net228 net455 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__mux2_1
XANTENNA__07007__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ net196 net1865 net410 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 net242 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 _04703_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
Xfanout262 _04696_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_4
XANTENNA__10052__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 _02712_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_2
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
XANTENNA__07715__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09841__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ net1158 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_198_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12822_ clknet_leaf_120_clk _00386_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12753_ clknet_leaf_110_clk _00317_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13660__Q net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11704_ _05525_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__xor2_2
XFILLER_0_84_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07494__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12684_ clknet_leaf_10_clk _00248_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11635_ _05482_ _05483_ _05474_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07246__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11566_ _05399_ _05408_ _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ clknet_leaf_36_clk _00869_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10517_ net2250 net257 net361 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10227__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ _05308_ net267 _05319_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07884__X _03011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13236_ clknet_leaf_45_clk _00800_ net1080 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ net150 net1778 net369 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
XANTENNA__08699__Y _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ clknet_leaf_20_clk _00731_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10379_ net429 net389 net385 net381 vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12118_ _05965_ _05977_ _05981_ _05984_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__nor4_1
X_13098_ clknet_leaf_38_clk _00662_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08221__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ _05890_ _05907_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_127_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06379__C top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10897__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06610_ top.DUT.register\[27\]\[28\] net778 net702 top.DUT.register\[29\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07590_ top.DUT.register\[22\]\[3\] net751 _01539_ top.DUT.register\[13\]\[3\] _02716_
+ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06541_ _01573_ net789 _01637_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__and3_4
XANTENNA__09703__B1_N net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06472_ net903 top.a1.instruction\[16\] top.a1.instruction\[19\] net900 vssd1 vssd1
+ vccd1 vccd1 _01599_ sky130_fd_sc_hd__and4_1
X_09260_ net894 _04293_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_173_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08211_ _02878_ net483 vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__or2_1
X_09191_ _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08142_ _02056_ net292 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07237__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08073_ _01713_ net291 _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10137__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07024_ top.DUT.register\[24\]\[11\] net551 net546 top.DUT.register\[5\]\[11\] _02150_
+ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08737__A2 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1023_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ net1258 net865 _01904_ net593 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a22o_1
XANTENNA__13745__Q top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 top.ramstore\[3\] vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_184_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 _01177_ vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold37 top.a1.row1\[18\] vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _03046_ _03048_ _03050_ _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__or4_2
Xhold48 top.a1.row1\[16\] vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold59 net122 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ top.DUT.register\[11\]\[18\] net642 net634 top.DUT.register\[19\]\[18\] _02983_
+ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout650_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ top.DUT.register\[17\]\[24\] net645 net621 top.DUT.register\[26\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a22o_1
XANTENNA__10600__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08277__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07788_ top.DUT.register\[25\]\[19\] net774 net687 top.DUT.register\[1\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09527_ net137 _04555_ _04561_ _04563_ net910 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__o221a_1
X_06739_ top.DUT.register\[26\]\[25\] net760 net686 top.DUT.register\[1\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_X clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09458_ net132 _04491_ _04497_ _04498_ top.i_ready vssd1 vssd1 vccd1 vccd1 _04499_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__07476__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08409_ net300 _03397_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__nand2_1
XANTENNA__06684__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net907 top.pc\[19\] _04433_ net896 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11420_ _05248_ _05254_ _05285_ _05251_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a22o_2
XFILLER_0_34_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07228__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11351_ _05182_ _05197_ top.a1.dataIn\[29\] vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__o21a_1
XANTENNA__10047__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06471__D top.a1.instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ net466 _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11282_ _05148_ _05150_ _05152_ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_95_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13021_ clknet_leaf_107_clk _00585_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10233_ _01601_ net466 _04929_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__nor3_4
XANTENNA__07864__B _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1020 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_4
X_10164_ net141 net1767 net416 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07400__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1013 net1019 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1024 net1029 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09138__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1035 net1038 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_2
Xfanout1046 net1050 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
Xfanout1057 net1060 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_2
X_10095_ net146 net1806 net418 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
Xfanout1068 net1084 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_2
XANTENNA__09689__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1079 net1084 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XFILLER_0_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12558__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ net1119 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XANTENNA__10510__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06496__A top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ clknet_leaf_116_clk _00369_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13785_ clknet_leaf_64_clk _01328_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08982__Y _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10997_ net1368 _05013_ net535 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12736_ clknet_leaf_46_clk _00300_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07467__A2 _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__B2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06675__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ clknet_leaf_47_clk _00231_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11618_ top.a1.dataIn\[11\] _05485_ _05486_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__or3_1
XANTENNA__07219__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12212__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ clknet_leaf_2_clk _00162_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08967__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ _05386_ _05417_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold507 top.DUT.register\[26\]\[0\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 top.DUT.register\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ clknet_leaf_22_clk _00783_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08760_ net888 top.pc\[22\] net537 _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a22o_1
X_13852__1117 vssd1 vssd1 vccd1 vccd1 _13852__1117/HI net1117 sky130_fd_sc_hd__conb_1
X_07711_ top.DUT.register\[29\]\[1\] net665 net614 top.DUT.register\[14\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a22o_1
X_08691_ net320 _03411_ _03543_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__a21bo_1
X_07642_ top.DUT.register\[27\]\[2\] net775 net678 top.DUT.register\[13\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a22o_1
XANTENNA__10420__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07573_ top.DUT.register\[29\]\[3\] net663 net651 top.DUT.register\[28\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09312_ _02380_ _04349_ _04353_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06524_ top.a1.instruction\[22\] top.a1.instruction\[23\] _01626_ vssd1 vssd1 vccd1
+ vccd1 _01651_ sky130_fd_sc_hd__o21a_1
XANTENNA__11714__D_N top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06666__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ top.pc\[11\] _02212_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__and2b_1
XFILLER_0_145_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06455_ _01579_ _01581_ _01576_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout329_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06386_ net792 _01511_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__nor2_4
X_09174_ _04228_ _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06418__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _03248_ _03251_ net276 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07091__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _03156_ _03160_ _03172_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__and3_4
XANTENNA__08413__X _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout698_A _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ top.DUT.register\[11\]\[11\] net758 net710 top.DUT.register\[9\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a22o_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__08132__Y _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__A_N top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07394__A1 top.a1.instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08958_ _02491_ net591 net1183 net865 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_90_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ top.DUT.register\[11\]\[16\] net756 net713 top.DUT.register\[30\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a22o_1
X_08889_ _01735_ net487 net470 _01736_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net218 net1666 net441 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XANTENNA__10330__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12850__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ net2195 net196 net351 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07449__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13570_ clknet_leaf_75_clk _01129_ net1088 vssd1 vssd1 vccd1 vccd1 top.a1.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08735__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ net1575 net222 net448 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06657__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ clknet_leaf_105_clk _00085_ net1001 vssd1 vssd1 vccd1 vccd1 top.pc\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12452_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[4\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08036__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12554__Q top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _05261_ _05263_ _05268_ _05270_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__o211ai_1
X_12383_ clknet_leaf_82_clk _00019_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11334_ _05189_ _05193_ top.a1.dataIn\[20\] vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07621__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ top.a1.row1\[122\] _05106_ _05120_ top.a1.row2\[42\] _05142_ vssd1 vssd1
+ vccd1 vccd1 _05143_ sky130_fd_sc_hd__a221o_1
XANTENNA__10505__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__Y _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13004_ clknet_leaf_10_clk _00568_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10216_ net179 net2022 net405 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ net1193 _05079_ _05085_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__a21o_1
XANTENNA__08582__B1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10147_ net195 net2129 net416 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
XANTENNA__09017__D _03652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__A2 _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10078_ net199 net2001 net419 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__mux2_1
XANTENNA__06497__Y _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10240__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06896__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ net72 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11860__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13768_ clknet_leaf_86_clk _01311_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ clknet_leaf_22_clk _00283_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ clknet_leaf_74_clk _01247_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06240_ net1280 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[16\] sky130_fd_sc_hd__and2_1
XANTENNA_wire499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07860__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06171_ wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold304 top.DUT.register\[18\]\[9\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold315 top.DUT.register\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 top.DUT.register\[24\]\[13\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 top.ramload\[25\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 top.DUT.register\[17\]\[12\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ net262 net2206 net433 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06820__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold359 top.DUT.register\[30\]\[16\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout806 net807 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_4
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_2
X_09861_ net169 net1594 net438 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__mux2_1
XANTENNA__08962__A2_N net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_4
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_0_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08812_ _03098_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_181_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09792_ top.pc\[19\] _04425_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__xnor2_1
Xhold1004 top.DUT.register\[2\]\[10\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06688__X _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1015 top.DUT.register\[21\]\[5\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 top.DUT.register\[6\]\[31\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1037 top.DUT.register\[2\]\[16\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net1317 net837 net816 _03848_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a22o_1
Xhold1048 top.DUT.register\[18\]\[17\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 top.DUT.register\[31\]\[7\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10150__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07679__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ net474 _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ top.DUT.register\[8\]\[2\] net568 net781 top.DUT.register\[31\]\[2\] _02751_
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_200_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10938__X _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A _04950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07556_ net319 _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_196_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06639__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ top.a1.instruction\[21\] net801 top.a1.instruction\[20\] vssd1 vssd1 vccd1
+ vccd1 _01634_ sky130_fd_sc_hd__and3b_2
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ top.DUT.register\[1\]\[5\] net655 net603 top.DUT.register\[18\]\[5\] _02613_
+ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_46_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07300__A1 top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ top.pc\[9\] top.pc\[10\] _04254_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__and3_1
X_06438_ top.a1.instruction\[6\] _01474_ top.a1.instruction\[2\] net905 vssd1 vssd1
+ vccd1 vccd1 _01565_ sky130_fd_sc_hd__nand4b_2
XANTENNA__07851__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13379__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09157_ _04214_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__nor2_1
X_06369_ top.a1.instruction\[17\] top.a1.instruction\[18\] net810 vssd1 vssd1 vccd1
+ vccd1 _01496_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ net287 _03225_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _01490_ _01571_ _01576_ _04147_ _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06811__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ _03127_ _03147_ _03164_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o211a_1
XANTENNA__10325__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 top.DUT.register\[8\]\[6\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12106__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 top.lcd.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08303__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold882 top.DUT.register\[25\]\[19\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net1264 net863 net827 top.ramstore\[1\] vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__a22o_1
Xhold893 top.DUT.register\[17\]\[21\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10001_ net251 net1823 net426 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06590__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10060__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ _05815_ _05820_ _05792_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06878__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10903_ net151 net1750 net441 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
X_11883_ _05736_ _05741_ net129 _05749_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13622_ clknet_leaf_75_clk net1277 net1088 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10834_ net2076 net147 net354 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__mux2_1
XANTENNA__08465__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ clknet_leaf_68_clk _01117_ net1104 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ net166 net1706 net376 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06493__B net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08037__Y _03164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12504_ clknet_leaf_61_clk _00071_ net1099 vssd1 vssd1 vccd1 vccd1 top.ramstore\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ clknet_leaf_11_clk _01048_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10696_ net190 net2252 net380 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
X_13851__1116 vssd1 vssd1 vccd1 vccd1 _13851__1116/HI net1116 sky130_fd_sc_hd__conb_1
XFILLER_0_82_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12435_ clknet_leaf_94_clk top.ru.next_FetchedData\[19\] net997 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09044__A1 _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07055__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12366_ _06148_ _06149_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ top.a1.dataIn\[19\] top.a1.dataIn\[18\] top.a1.dataIn\[17\] top.a1.dataIn\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10235__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] top.lcd.cnt_500hz\[6\] _01438_
+ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_73_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248_ top.a1.row2\[32\] _05107_ _05122_ _05127_ _05104_ vssd1 vssd1 vccd1 vccd1
+ _05128_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ top.a1.dataInTemp\[11\] top.a1.data\[11\] net799 vssd1 vssd1 vccd1 vccd1
+ _05077_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06581__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12459__Q top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07410_ top.DUT.register\[17\]\[7\] net644 net564 top.DUT.register\[4\]\[7\] _02526_
+ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a221o_1
X_08390_ _03494_ _03495_ net283 vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07341_ _02463_ _02465_ _02467_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07294__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ net807 _02398_ _01624_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07833__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _03658_ _03586_ _03632_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and3b_1
XFILLER_0_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06223_ net2012 _01404_ top.Wen wb.curr_state\[2\] net918 vssd1 vssd1 vccd1 vccd1
+ _00016_ sky130_fd_sc_hd__a32o_1
XANTENNA__09035__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06154_ top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XANTENNA__07046__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 _01184_ vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09586__A2 _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold112 top.DUT.register\[4\]\[10\] vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold123 top.a1.row1\[12\] vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold134 top.ramaddr\[7\] vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 top.DUT.register\[11\]\[3\] vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10145__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 top.a1.row2\[12\] vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 top.a1.row2\[9\] vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09934__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ net835 _04604_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__o21ba_1
Xhold178 top.a1.row1\[106\] vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _01668_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_74_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold189 top.a1.row1\[105\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _01666_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
Xfanout625 _01662_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _01652_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_2
Xfanout647 _01642_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_8
X_09844_ net833 _04506_ _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__o21bai_1
XANTENNA__07962__B _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 _01639_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08010__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _01554_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_8
X_09775_ _04769_ _04772_ _04778_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__o21ai_1
X_06987_ top.DUT.register\[11\]\[20\] net642 net628 top.DUT.register\[9\]\[20\] _02113_
+ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a221o_1
XANTENNA__13753__Q top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout563_A _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06572__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ net888 top.pc\[20\] net537 _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a22o_1
XANTENNA__08849__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10656__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08657_ _03342_ _03542_ _03582_ net270 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout730_A _01523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout828_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ top.a1.instruction\[9\] _01477_ _01620_ top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 _02735_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_194_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _03646_ _03700_ net278 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07539_ top.DUT.register\[11\]\[4\] net757 net687 top.DUT.register\[1\]\[4\] _02665_
+ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a221o_1
XFILLER_0_181_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_10__f_clk_X clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ net257 net1637 net357 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__mux2_1
XANTENNA__07285__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ _04263_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__nand2_1
XANTENNA__09026__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ net148 net2269 net365 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__mux2_1
X_12220_ net1181 _06053_ net589 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
X_12151_ _06005_ _06015_ _06014_ _06011_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10055__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ net914 net1347 net854 _05037_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__a31o_1
XFILLER_0_208_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12082_ top.a1.dataIn\[3\] _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__and2b_1
Xhold690 top.DUT.register\[16\]\[3\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
X_11033_ net12 net831 net830 top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__a22o_1
XANTENNA__08001__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__A _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__A2 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12984_ clknet_leaf_109_clk _00548_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08984__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11935_ _05776_ _05782_ _05791_ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a31o_1
XFILLER_0_200_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11866_ _05728_ _05734_ _05721_ _05724_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_156_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13605_ clknet_leaf_95_clk _01164_ net990 vssd1 vssd1 vccd1 vccd1 top.ramload\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_205_Right_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817_ net1507 net202 net355 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11797_ _05572_ _05605_ _05628_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08208__B _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ clknet_leaf_49_clk _01100_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10748_ net231 net1771 net374 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__mux2_1
XANTENNA__07815__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13467_ clknet_leaf_58_clk _01031_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ net253 net2169 net379 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07028__B1 _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12418_ clknet_leaf_96_clk top.ru.next_FetchedData\[2\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_132_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13398_ clknet_leaf_2_clk _00962_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07579__A1 top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__B1 _03875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12349_ _06137_ _06138_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__nor2_1
XANTENNA__12891__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06910_ _02035_ _02036_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__nor2_2
X_07890_ top.DUT.register\[4\]\[17\] net564 net548 top.DUT.register\[24\]\[17\] _03016_
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a221o_1
XANTENNA__07200__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06841_ top.DUT.register\[30\]\[23\] net615 net540 top.DUT.register\[22\]\[23\] _01967_
+ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06554__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ net910 net897 _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_90_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06772_ top.DUT.register\[1\]\[25\] net656 net620 top.DUT.register\[26\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08511_ net522 _03626_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_160_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09491_ _04527_ _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08442_ _03228_ _03249_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08373_ _03365_ _03369_ net298 vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_176_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout144_A _04908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07324_ top.DUT.register\[27\]\[8\] net775 net731 top.DUT.register\[19\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07267__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09929__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07806__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07255_ top.DUT.register\[17\]\[14\] net645 net547 top.DUT.register\[5\]\[14\] _02381_
+ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout311_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07019__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06206_ top.busy_o top.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 top.ru.next_iready sky130_fd_sc_hd__and2b_1
XFILLER_0_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07186_ top.DUT.register\[2\]\[13\] net661 net646 top.DUT.register\[17\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13748__Q top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07973__A _01865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _04941_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_8
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XANTENNA__08519__B1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout778_A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _04925_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06793__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 _04918_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10603__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 _04965_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 _04936_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_4
Xfanout466 _04676_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_8
X_09827_ _04476_ net526 net332 top.a1.dataIn\[22\] net334 vssd1 vssd1 vccd1 vccd1
+ _04828_ sky130_fd_sc_hd__a221o_1
Xfanout477 _03330_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_129_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout945_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06545__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850__1115 vssd1 vssd1 vccd1 vccd1 _13850__1115/HI net1115 sky130_fd_sc_hd__conb_1
X_09758_ _01567_ _04372_ _04379_ net527 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_87_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _03780_ _03815_ _02949_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a21o_1
XFILLER_0_201_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _03490_ net341 net338 _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__o211a_2
XFILLER_0_139_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12591__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ _01395_ _05559_ _05528_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11651_ _05494_ _05498_ _05519_ _05497_ _05481_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ net175 net2190 net385 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09798__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11582_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13321_ clknet_leaf_4_clk _00885_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10533_ net1457 net203 net363 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__mux2_1
XANTENNA__08470__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_clk_X clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_40_clk _00816_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10464_ net229 net1756 net370 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__mux2_1
XANTENNA__08044__A _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13658__Q net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12203_ _05922_ _04976_ net847 top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 _01288_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_114_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13183_ clknet_leaf_114_clk _00747_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ net199 net1827 net329 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__mux2_1
XANTENNA__07430__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ _05989_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_209_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08731__A2_N net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06784__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ _05918_ _05920_ _05933_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08050__Y _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ net24 net832 net830 net1890 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__a22o_1
XANTENNA__09722__A2 _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08930__B1 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__B _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12967_ clknet_leaf_27_clk _00531_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13437__RESET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _05754_ _05763_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07497__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12898_ clknet_leaf_42_clk _00462_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11849_ _05688_ _05713_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or3_1
XANTENNA__09238__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07249__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07777__B _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ clknet_leaf_22_clk _01083_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload10 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload21 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload21/X sky130_fd_sc_hd__clkbuf_4
X_07040_ top.DUT.register\[22\]\[10\] net752 net705 top.DUT.register\[15\]\[10\] _02166_
+ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload32 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__inv_6
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload43 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_58_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12472__Q top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload54 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__clkinv_4
Xclkload65 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__clkinv_8
Xclkload76 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_4
Xclkload87 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload87/X sky130_fd_sc_hd__clkbuf_4
Xclkload98 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07421__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08991_ _03557_ _03592_ _03614_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and4_1
XANTENNA__06775__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07972__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ top.DUT.register\[28\]\[16\] net652 net567 top.DUT.register\[4\]\[16\] _03057_
+ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a221o_1
XANTENNA__10423__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07873_ top.DUT.register\[12\]\[17\] net580 net751 top.DUT.register\[22\]\[17\] _02994_
+ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09612_ top.a1.state\[1\] _04639_ _04642_ _04631_ vssd1 vssd1 vccd1 vccd1 _00114_
+ sky130_fd_sc_hd__o22a_1
X_06824_ _01929_ _01949_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__and2_1
XANTENNA__07017__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09543_ _01755_ _04577_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__nor2_1
X_06755_ top.DUT.register\[19\]\[25\] net734 net718 top.DUT.register\[2\]\[25\] _01876_
+ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__A1 top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08886__A1_N net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07488__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net132 _04504_ _04505_ _04513_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09232__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06686_ top.DUT.register\[29\]\[27\] net664 net619 top.DUT.register\[26\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a22o_1
XANTENNA__08129__A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__B net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ net311 net490 vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__or2_2
XFILLER_0_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _03341_ _03477_ net307 vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__X _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload4/X sky130_fd_sc_hd__clkbuf_2
X_07307_ top.DUT.register\[13\]\[9\] net648 net636 top.DUT.register\[16\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ net284 _03410_ _03407_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07238_ top.DUT.register\[15\]\[14\] net706 _02362_ _02364_ vssd1 vssd1 vccd1 vccd1
+ _02365_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07169_ top.DUT.register\[17\]\[13\] net724 net676 top.DUT.register\[18\]\[13\] _02295_
+ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08799__A _01909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ net200 net1482 net411 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10333__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _04775_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09165__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout252 _04703_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_1
Xfanout263 net266 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_4
XFILLER_0_199_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout285 _02712_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
Xfanout296 _02810_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlymetal6s2s_1
X_13870_ net1157 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_198_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12821_ clknet_leaf_6_clk _00385_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09468__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12752_ clknet_leaf_121_clk _00316_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07479__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11275__A1 top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08676__C1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ _05529_ _05531_ _05559_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12557__Q top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12683_ clknet_leaf_30_clk _00247_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11634_ _05488_ _05489_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08979__B1 _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11565_ _05388_ _05396_ _05397_ net250 _05394_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a41o_1
XANTENNA__10508__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13304_ clknet_leaf_112_clk _00868_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10516_ net1578 net261 net361 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__mux2_1
X_11496_ _05365_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13235_ clknet_leaf_4_clk _00799_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ _04676_ _04680_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__nand2_8
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07403__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ clknet_leaf_116_clk _00730_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ net450 net377 _04951_ net373 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__and4b_1
X_12117_ _05977_ _05981_ _05984_ _05986_ _05978_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__o32a_1
XANTENNA__07954__B2 _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ clknet_leaf_3_clk _00661_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08221__B net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ _05913_ _05916_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08903__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07182__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09459__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13271__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06540_ _01640_ _01645_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__nor2_4
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06471_ top.a1.instruction\[25\] top.a1.instruction\[26\] top.a1.instruction\[27\]
+ top.a1.instruction\[28\] vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__and4_1
XFILLER_0_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08210_ _02881_ _03333_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__nand2_1
XANTENNA__07890__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09190_ _04228_ _04229_ _04230_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06692__A _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ _03265_ _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__nand2_1
XANTENNA__10418__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08072_ _01755_ net294 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__nand2_1
XANTENNA__07642__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07023_ top.DUT.register\[8\]\[11\] net570 net618 top.DUT.register\[30\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08412__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10153__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ net515 net592 net1188 net868 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__a2bb2o_1
X_13864__1125 vssd1 vssd1 vccd1 vccd1 _13864__1125/HI net1125 sky130_fd_sc_hd__conb_1
XANTENNA_fanout1016_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08131__B _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 _01170_ vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09942__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold27 top.lcd.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ top.DUT.register\[31\]\[16\] net744 net690 top.DUT.register\[3\]\[16\] _03051_
+ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a221o_1
Xhold38 top.ramstore\[28\] vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 top.a1.row1\[17\] vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ top.DUT.register\[3\]\[18\] net788 _02982_ vssd1 vssd1 vccd1 vccd1 _02983_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07173__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ top.DUT.register\[21\]\[24\] net575 net625 top.DUT.register\[25\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07787_ top.DUT.register\[31\]\[19\] net745 net695 top.DUT.register\[21\]\[19\] _02913_
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout643_A _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06920__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ _01618_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06738_ _01861_ _01863_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__nor2_2
XFILLER_0_183_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ _04492_ _04496_ _01619_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a21o_1
XFILLER_0_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06669_ _01784_ _01785_ _01794_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__or4_4
XANTENNA__09897__B _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ net301 _03400_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12206__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06185__A_N top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07881__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ net139 _04415_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08339_ _03458_ _03461_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__or2_2
XFILLER_0_191_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10328__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11013__A top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _05217_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06987__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ _04679_ _04937_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11281_ net891 top.a1.row1\[115\] _05105_ _05156_ _05157_ vssd1 vssd1 vccd1 vccd1
+ _05158_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_111_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09386__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ clknet_leaf_17_clk _00584_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09418__A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10232_ net141 net2024 net407 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__mux2_1
XANTENNA__06739__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ net144 net2329 net414 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08041__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1014 net1016 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 net1029 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09852__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__X _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1036 net1038 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
Xfanout1047 net1050 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_2
XANTENNA_input37_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09689__A1 _03490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ net152 net1608 net419 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
Xfanout1058 net1060 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
Xfanout1069 net1076 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ net1118 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_186_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06911__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06496__B _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ clknet_leaf_40_clk _00368_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11248__A1 top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ clknet_leaf_64_clk _01327_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10996_ top.a1.dataIn\[7\] net848 net843 _05012_ vssd1 vssd1 vccd1 vccd1 _05013_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ clknet_leaf_115_clk _00299_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07872__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ clknet_leaf_18_clk _00230_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08056__X _03183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11617_ _05485_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__or2_1
XANTENNA__10238__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ clknet_leaf_6_clk _00161_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09613__A1 _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ _05382_ _05386_ net250 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__or3b_1
XFILLER_0_107_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06978__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 top.DUT.register\[5\]\[23\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold519 top.DUT.register\[24\]\[16\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ _05342_ _05343_ _05347_ _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__o31a_2
XANTENNA__08503__Y _03619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13218_ clknet_leaf_42_clk _00782_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08232__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13149_ clknet_leaf_107_clk _00713_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ top.DUT.register\[15\]\[1\] _01655_ net784 top.DUT.register\[31\]\[1\] _02836_
+ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a221o_1
X_08690_ _02951_ _03085_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10701__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07155__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ top.DUT.register\[19\]\[2\] net731 net689 top.DUT.register\[3\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07572_ top.DUT.register\[20\]\[3\] net576 net635 top.DUT.register\[16\]\[3\] _02698_
+ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09311_ _04357_ _04358_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__xor2_1
XANTENNA__09301__B1 _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06523_ _01590_ _01628_ net789 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_157_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10937__A _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _04293_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06454_ _01479_ _01580_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nand2_2
XANTENNA__07863__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09173_ _04229_ _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nand2_1
X_06385_ net791 _01511_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__nor2_4
XANTENNA__10148__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ _03249_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09937__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07615__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06969__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _03156_ _03160_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07006_ top.DUT.register\[28\]\[11\] net587 net694 top.DUT.register\[21\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
XANTENNA__08142__A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09672__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ net1267 net865 _02540_ net593 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout760_A _01510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _03033_ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__nor2_2
X_08888_ _03675_ _03771_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nor2_1
X_07839_ top.DUT.register\[12\]\[18\] net583 net710 top.DUT.register\[9\]\[18\] _02965_
+ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a221o_1
XFILLER_0_196_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ net2108 net201 net352 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09509_ _04544_ _04545_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__xor2_1
X_10781_ net1669 net223 net445 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ clknet_leaf_80_clk _00084_ net1002 vssd1 vssd1 vccd1 vccd1 top.pc\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07854__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08317__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[3\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[3\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__10058__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ _05265_ _05268_ _05270_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12382_ clknet_leaf_88_clk _00018_ net1005 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ top.a1.dataIn\[23\] _05189_ _05191_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08323__Y _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ top.a1.row1\[10\] _05108_ _05112_ top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1
+ _05142_ sky130_fd_sc_hd__a22o_1
X_13003_ clknet_leaf_31_clk _00567_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10215_ net195 net2207 net407 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__mux2_1
X_11195_ net851 _05071_ _05078_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and3_1
XANTENNA__07385__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ net202 net1597 net416 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06593__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10521__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ net208 net1776 net419 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08334__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07137__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload2_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13836_ clknet_leaf_68_clk _01377_ net1106 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13767_ clknet_leaf_86_clk _01310_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10979_ top.a1.halfData\[2\] _04991_ _05000_ net843 vssd1 vssd1 vccd1 vccd1 _05001_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07845__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ clknet_leaf_116_clk _00282_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13863__1124 vssd1 vssd1 vccd1 vccd1 _13863__1124/HI net1124 sky130_fd_sc_hd__conb_1
XFILLER_0_45_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13698_ clknet_leaf_73_clk _01246_ net1091 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12649_ clknet_leaf_2_clk _00213_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09757__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06170_ net1 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13300__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold305 top.DUT.register\[26\]\[14\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12195__A2_N _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 top.DUT.register\[6\]\[1\] vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold327 top.DUT.register\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 top.DUT.register\[23\]\[9\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 top.DUT.register\[14\]\[8\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout807 _01563_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
X_09860_ net337 _04851_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and3_4
Xfanout818 _03264_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_2
Xfanout829 _05026_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_4
XANTENNA__07376__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ _01909_ _03097_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__nand2_1
X_09791_ net214 top.DUT.register\[1\]\[18\] net440 vssd1 vssd1 vccd1 vccd1 _00140_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06584__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 top.DUT.register\[30\]\[14\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 top.DUT.register\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 top.DUT.register\[2\]\[7\] vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ net888 top.pc\[21\] net537 _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a22o_1
Xhold1038 top.DUT.register\[12\]\[6\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10431__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1049 top.DUT.register\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08325__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08673_ _03780_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_163_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout174_A _04850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07624_ top.DUT.register\[19\]\[2\] net631 net779 top.DUT.register\[15\]\[2\] _02741_
+ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07555_ _02674_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_37_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout341_A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1083_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _04681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06506_ _01629_ _01632_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nor2_8
XANTENNA__07836__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07486_ top.DUT.register\[13\]\[5\] net647 net635 top.DUT.register\[16\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09225_ net909 top.pc\[9\] _04279_ net897 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_101_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06437_ top.a1.instruction\[6\] _01474_ top.a1.instruction\[2\] net905 vssd1 vssd1
+ vccd1 vccd1 _01564_ sky130_fd_sc_hd__and4b_1
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_A _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09156_ top.pc\[5\] _02641_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__and2_1
X_06368_ _01476_ _01494_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08107_ net276 _03169_ _03226_ net300 vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ net833 _02201_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and3_1
XANTENNA__10606__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06299_ net2298 _01445_ _01446_ net892 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__a22oi_4
Xclkbuf_leaf_110_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ _03160_ _03156_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold850 top.DUT.register\[4\]\[21\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 top.DUT.register\[20\]\[12\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08303__C _03426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08013__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 top.DUT.register\[21\]\[21\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 top.DUT.register\[2\]\[15\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 top.DUT.register\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ net255 net2160 net425 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_110_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06575__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ net2255 net160 net429 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
XANTENNA__10341__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _05815_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_106_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10902_ _01601_ net465 _04937_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__or3b_4
XFILLER_0_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11882_ top.a1.dataIn\[5\] _05750_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__xor2_2
XANTENNA__08469__A2_N net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__A top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13621_ clknet_leaf_75_clk net1211 net1090 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
X_10833_ net1510 net153 net355 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__mux2_1
XANTENNA__08619__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07827__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13552_ clknet_leaf_72_clk _01116_ net1095 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_10764_ net169 net1885 net374 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08047__A _03164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ clknet_leaf_45_clk _00070_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramstore\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13483_ clknet_leaf_31_clk _01047_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net194 net1543 net379 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ clknet_leaf_92_clk top.ru.next_FetchedData\[18\] net1000 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[18\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_43_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12365_ net1356 _06146_ net796 vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10516__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11316_ top.a1.dataIn\[31\] top.a1.dataIn\[25\] top.a1.dataIn\[24\] top.a1.dataIn\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nand4_1
X_12296_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] _01438_ top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ top.a1.row2\[16\] _05118_ _05124_ _05126_ vssd1 vssd1 vccd1 vccd1 _05127_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08004__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__A1 _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output68_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net1334 net532 net525 _05076_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a22o_1
XANTENNA__08510__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10251__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net1395 net142 net460 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10114__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07413__X _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ clknet_leaf_67_clk _01360_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09807__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07340_ top.DUT.register\[10\]\[8\] net727 net700 top.DUT.register\[29\]\[8\] _02466_
+ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07818__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12475__Q top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07271_ _02382_ _02395_ _02396_ _02397_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__or4_2
XFILLER_0_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09010_ _03412_ _03546_ _03566_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06222_ wb.curr_state\[0\] top.Ren _01405_ net2120 net918 vssd1 vssd1 vccd1 vccd1
+ _00015_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09035__A2 _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06153_ net2125 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10426__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 top.ramaddr\[18\] vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 top.ramaddr\[16\] vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__B _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 net86 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 top.DUT.register\[31\]\[25\] vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 top.ramaddr\[11\] vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 top.ramaddr\[21\] vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 top.ramaddr\[17\] vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _04605_ net526 net333 top.a1.dataIn\[30\] net335 vssd1 vssd1 vccd1 vccd1
+ _04905_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_74_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold179 top.a1.row1\[107\] vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout604 _01668_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08546__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout615 _01664_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07349__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout626 _01662_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _04508_ net526 net332 top.a1.dataIn\[24\] net334 vssd1 vssd1 vccd1 vccd1
+ _04842_ sky130_fd_sc_hd__a221o_1
Xfanout637 _01652_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06557__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 _01642_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_4
XANTENNA_fanout291_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _01638_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout389_A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10161__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06986_ top.DUT.register\[15\]\[20\] net780 _02100_ _02112_ vssd1 vssd1 vccd1 vccd1
+ _02113_ sky130_fd_sc_hd__a211o_1
X_09774_ _04769_ _04772_ _04777_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09950__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07036__A _02142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ _03821_ _03829_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_198_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout556_A _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _03680_ _03765_ net307 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07521__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ top.a1.instruction\[23\] _01617_ _01621_ top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
X_08587_ _03239_ _03243_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nand2_1
XANTENNA__09259__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A _01527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07538_ top.DUT.register\[31\]\[4\] net745 net709 top.DUT.register\[9\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07809__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ top.DUT.register\[8\]\[5\] net739 net716 top.DUT.register\[2\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ net500 _02471_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__nand2_1
X_10480_ _04676_ _04917_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__nand2_8
XFILLER_0_134_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09026__A2 _03483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ top.pc\[4\] _04182_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07588__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ net41 net858 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__and2_1
X_12081_ _05912_ _05946_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__xnor2_2
Xhold680 top.DUT.register\[20\]\[8\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 top.DUT.register\[31\]\[10\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net11 net831 net830 net1386 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__a22o_1
XANTENNA__11136__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__A top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862__1123 vssd1 vssd1 vccd1 vccd1 _13862__1123/HI net1123 sky130_fd_sc_hd__conb_1
XANTENNA__10071__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__B _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__A2 _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12983_ clknet_leaf_106_clk _00547_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08984__B _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ _05779_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09161__A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ _05721_ _05724_ _05728_ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06720__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13604_ clknet_leaf_95_clk _01163_ net988 vssd1 vssd1 vccd1 vccd1 top.ramload\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ net1444 net208 net355 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11796_ _05664_ _05610_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__and2b_1
XANTENNA__08961__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ clknet_leaf_111_clk _01099_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10747_ net237 top.DUT.register\[26\]\[8\] net373 vssd1 vssd1 vccd1 vccd1 _00930_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09670__C1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10678_ net255 net1821 net377 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__mux2_1
X_13466_ clknet_leaf_18_clk _01030_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08505__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12417_ clknet_leaf_96_clk top.ru.next_FetchedData\[1\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_180_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10246__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ clknet_leaf_7_clk _00961_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07579__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__A1 _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08776__B2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ _01403_ _06136_ net796 vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06787__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_206_Left_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12279_ top.lcd.cnt_20ms\[16\] top.lcd.cnt_20ms\[15\] _06092_ vssd1 vssd1 vccd1 vccd1
+ _06096_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08511__Y _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06840_ top.DUT.register\[6\]\[23\] net556 net631 top.DUT.register\[19\]\[23\] _01966_
+ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a221o_1
XANTENNA__07127__Y _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06771_ top.DUT.register\[28\]\[25\] net652 net549 top.DUT.register\[24\]\[25\] _01897_
+ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a221o_1
X_08510_ net317 _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_160_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ _04502_ _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__and2_1
X_08441_ net316 _03559_ _03558_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06711__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08372_ _02890_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07323_ _02448_ _02449_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11063__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07254_ top.DUT.register\[20\]\[14\] net578 net665 top.DUT.register\[29\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06205_ top.ru.state\[4\] net2030 top.busy_o vssd1 vssd1 vccd1 vccd1 top.ru.next_dready
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07185_ top.DUT.register\[8\]\[13\] net570 net550 top.DUT.register\[24\]\[13\] _02311_
+ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a221o_1
XANTENNA__10156__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1046_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09945__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06778__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _04939_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_8
Xfanout412 _04933_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09716__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 _04925_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_6
Xfanout434 _04918_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
Xfanout445 _04950_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_8
Xfanout456 net458 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_6
X_09826_ _04823_ _04825_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout478 _03257_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_4
Xfanout489 _03178_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09680__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07742__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09757_ net179 net1981 net438 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06969_ top.DUT.register\[1\]\[20\] net688 net679 top.DUT.register\[13\]\[20\] _02095_
+ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _02950_ _02991_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__nor2_1
X_09688_ net344 _04705_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__or2_1
X_08639_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11650_ _05494_ _05498_ _05519_ _05497_ _05481_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12886__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ net183 net1965 net387 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
X_11581_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10532_ net1759 net211 net364 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ clknet_leaf_31_clk _00884_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ clknet_leaf_50_clk _00815_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10463_ net180 net1888 net369 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10066__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _05946_ _04976_ net847 net2327 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_114_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09708__X _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ clknet_leaf_14_clk _00746_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10394_ net209 top.DUT.register\[15\]\[12\] net330 vssd1 vssd1 vccd1 vccd1 _00582_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06769__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _05998_ _06000_ _05994_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09707__B1 _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _05893_ _05900_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__or2_1
XANTENNA__08060__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ net13 net832 _05024_ net2102 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__a22o_1
XANTENNA__07194__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 net996 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07733__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06941__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12966_ clknet_leaf_19_clk _00530_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11917_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12897_ clknet_leaf_27_clk _00461_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11848_ _05681_ _05685_ _05686_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11779_ _05647_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13518_ clknet_leaf_111_clk _01082_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload11 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_153_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13449_ clknet_leaf_3_clk _01013_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload22 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_140_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload33 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload44 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_58_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload55 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload66 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinv_4
Xclkload77 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_6
Xclkload88 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_4
Xclkload99 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload99/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10704__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ _03421_ _03488_ _03518_ _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_71_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07941_ _03060_ _03062_ _03064_ _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07872_ top.DUT.register\[14\]\[17\] net720 net667 top.DUT.register\[5\]\[17\] _02998_
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07185__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ net893 _04639_ _04641_ _04642_ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__o22a_1
X_06823_ _01929_ _01949_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06932__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09542_ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__inv_2
X_06754_ top.DUT.register\[9\]\[25\] net709 net680 top.DUT.register\[13\]\[25\] _01878_
+ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09473_ net819 _04511_ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__or3_1
X_06685_ _01805_ _01807_ _01809_ _01811_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__or4_1
XANTENNA__08685__B1 _03793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_A _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08424_ _03542_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _03422_ _03476_ net281 vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout421_A _04925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13147__RESET_B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ top.DUT.register\[12\]\[9\] net608 net604 top.DUT.register\[18\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a22o_1
Xclkload5 clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_8
X_13861__1122 vssd1 vssd1 vccd1 vccd1 _13861__1122/HI net1122 sky130_fd_sc_hd__conb_1
X_08286_ net299 _03408_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_22_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06999__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07237_ top.DUT.register\[14\]\[14\] net723 net718 top.DUT.register\[2\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07168_ top.DUT.register\[26\]\[13\] net761 net706 top.DUT.register\[15\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XANTENNA__08432__X _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10614__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ top.DUT.register\[16\]\[10\] net636 net630 top.DUT.register\[9\]\[10\] _02213_
+ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a221o_1
Xfanout220 _04732_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_1
Xfanout231 _04726_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 _04715_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 _04703_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07176__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _03188_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
XANTENNA__08912__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07715__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09809_ net193 net2324 net440 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__mux2_1
Xfanout297 _02810_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ clknet_leaf_46_clk _00384_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12751_ clknet_leaf_21_clk _00315_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10483__A0 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11702_ _05550_ _05566_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12682_ clknet_leaf_38_clk _00246_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11633_ _05501_ _05502_ _05470_ _05484_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08979__B2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ _05424_ _05430_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__or2_1
XANTENNA__10786__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07100__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ clknet_leaf_106_clk _00867_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10515_ net1373 net263 net363 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__mux2_1
X_11495_ _05305_ _05355_ _05354_ _05307_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_150_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13234_ clknet_leaf_48_clk _00798_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10446_ net140 top.DUT.register\[16\]\[31\] net325 vssd1 vssd1 vccd1 vccd1 _00633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10377_ net466 _04934_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__nand2_8
XANTENNA__10524__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13165_ clknet_leaf_25_clk _00729_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12901__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12116_ _05967_ _05975_ _05966_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a21oi_1
X_13096_ clknet_leaf_34_clk _00660_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12047_ _05848_ _05903_ _05912_ _05915_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__and4_1
XANTENNA__08903__A1 _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output50_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06914__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12040__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13658__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ clknet_leaf_5_clk _00513_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06470_ top.a1.instruction\[10\] top.a1.instruction\[11\] _01508_ _01595_ vssd1 vssd1
+ vccd1 vccd1 _01597_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13240__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08140_ _01991_ net292 vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12483__Q top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload100 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__inv_12
X_08071_ net298 _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or2_1
XANTENNA__11103__B net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07022_ top.DUT.register\[20\]\[11\] net579 net562 top.DUT.register\[23\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Left_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10434__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ net1934 net866 _01972_ _04043_ vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 top.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 top.ramstore\[24\] vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ top.DUT.register\[8\]\[16\] net740 net673 top.DUT.register\[16\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a22o_1
Xhold39 _01195_ vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ top.DUT.register\[31\]\[18\] net784 net780 top.DUT.register\[15\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a22o_1
XANTENNA__06905__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A _04958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A _03339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09243__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ top.DUT.register\[1\]\[24\] net657 net617 top.DUT.register\[30\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_166_Left_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07786_ top.DUT.register\[6\]\[19\] net765 net761 top.DUT.register\[26\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_203_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ _04560_ _04559_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__nand2b_1
X_06737_ _01863_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout636_A _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ _04492_ _04496_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nor2_1
X_06668_ top.DUT.register\[18\]\[27\] net674 net671 top.DUT.register\[16\]\[27\] _01779_
+ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a221o_1
XANTENNA__07330__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _03395_ _03404_ net301 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06684__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07881__B2 top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ net135 _04421_ _04430_ _04431_ net907 vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__o221a_1
XANTENNA__12206__B2 top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06599_ _01717_ _01719_ _01721_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ net478 _03448_ _03449_ _03334_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ net280 _03277_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07633__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_175_Left_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10300_ net1665 net140 net403 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ top.a1.row2\[43\] _05120_ _05100_ _01444_ vssd1 vssd1 vccd1 vccd1 _05157_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_111_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10231_ net144 net1357 net406 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10344__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ net153 net1794 net415 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
Xfanout1004 net1020 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_7_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09138__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_2
Xfanout1026 net1029 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_2
X_10093_ net158 net2259 net420 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_2
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
Xfanout1059 net1060 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09689__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__X _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_184_Left_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ net1117 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ clknet_leaf_22_clk _00367_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13783_ clknet_leaf_64_clk _01326_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10995_ top.a1.data\[3\] top.a1.dataInTemp\[7\] net797 vssd1 vssd1 vccd1 vccd1 _05012_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12734_ clknet_leaf_14_clk _00298_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06675__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12665_ clknet_leaf_37_clk _00229_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10519__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11204__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11616_ top.a1.dataIn\[12\] _05482_ _05483_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__and3_1
XFILLER_0_182_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ clknet_leaf_60_clk _00160_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08870__A1_N net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11547_ _05381_ _05407_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold509 top.DUT.register\[27\]\[10\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xwire495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_8
X_11478_ _05328_ _05343_ _05329_ _05325_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09377__A1 _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ clknet_leaf_27_clk _00781_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10254__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ net197 net2095 net325 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13148_ clknet_leaf_54_clk _00712_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13079_ clknet_leaf_17_clk _00643_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_183_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07416__X _02543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07640_ top.DUT.register\[17\]\[2\] net726 net696 top.DUT.register\[23\]\[2\] _02766_
+ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a221o_1
XANTENNA__12478__Q top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ top.DUT.register\[13\]\[3\] net647 net643 top.DUT.register\[17\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06522_ _01629_ _01645_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__nor2_1
X_09310_ _04357_ _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_24_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07312__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06453_ net903 net901 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__nand2_1
X_09241_ top.pc\[11\] _04280_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06666__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12947__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09172_ _02612_ top.pc\[6\] vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__nand2b_1
X_06384_ net810 _01505_ _01508_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__nand3_2
XFILLER_0_113_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08123_ net503 net289 vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__nand2_1
XANTENNA__06418__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ _03169_ _03177_ net483 _03170_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07091__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ top.DUT.register\[6\]\[11\] net766 net725 top.DUT.register\[17\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10164__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07379__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout586_A _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ net1195 net869 _02585_ net594 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_205_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07907_ _03012_ _03032_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__nor2_1
X_08887_ net318 _03683_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a21o_2
XANTENNA_fanout753_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09540__A1 top.a1.instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ top.DUT.register\[15\]\[18\] net707 net703 top.DUT.register\[29\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _02279_ _02404_ _02450_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_36_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09508_ _04545_ _04544_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10780_ net1970 net233 net446 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07303__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ net136 _04470_ _04479_ _04480_ net906 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06657__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10339__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08054__A2_N _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[2\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_97_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11401_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12381_ clknet_leaf_71_clk net1165 net1093 vssd1 vssd1 vccd1 vccd1 top.edg2.flip2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _05191_ _05194_ top.a1.dataIn\[23\] vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10074__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ net880 _05103_ _05113_ top.a1.row2\[26\] _05140_ vssd1 vssd1 vccd1 vccd1
+ _05141_ sky130_fd_sc_hd__a221o_1
X_13002_ clknet_leaf_34_clk _00566_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07909__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ net200 net2290 net407 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09716__X _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11194_ net1243 net530 _05084_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__a21o_1
XANTENNA__08620__X _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__A2 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ net207 net2116 net413 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_192_Left_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10802__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07790__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ net222 top.DUT.register\[6\]\[11\] net419 vssd1 vssd1 vccd1 vccd1 _00293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08334__A2 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07542__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13835_ clknet_leaf_68_clk _01376_ net1106 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06896__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_48_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13766_ clknet_leaf_85_clk _01309_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ top.a1.dataInTemp\[2\] net799 vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ clknet_leaf_32_clk _00281_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10249__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ clknet_leaf_73_clk _01245_ net1091 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12648_ clknet_leaf_35_clk _00212_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12579_ clknet_leaf_50_clk _00143_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 top.DUT.register\[13\]\[27\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 top.DUT.register\[31\]\[16\] vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 top.DUT.register\[27\]\[2\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold339 top.DUT.register\[20\]\[1\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06820__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
Xfanout819 _01588_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_4
X_08810_ net275 net519 _03296_ _03908_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o311a_1
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10712__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _03794_ net340 net336 _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__o211a_4
XANTENNA__13683__SET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 top.DUT.register\[28\]\[1\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 top.DUT.register\[17\]\[9\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net474 _03835_ _03846_ net471 _03845_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__o221ai_4
XPHY_EDGE_ROW_183_Right_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1028 top.pad.keyCode\[2\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 top.lcd.currentState\[2\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
X_08672_ _02993_ _03779_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_163_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09361__X _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ top.DUT.register\[2\]\[2\] net659 net619 top.DUT.register\[26\]\[2\] _02749_
+ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a221o_1
XANTENNA__09802__A top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10948__A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout167_A _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ _02676_ _02678_ _02680_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__or3_1
XANTENNA__09521__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08418__A _03537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07322__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06505_ top.a1.instruction\[20\] top.a1.instruction\[21\] net900 _01626_ vssd1 vssd1
+ vccd1 vccd1 _01632_ sky130_fd_sc_hd__or4bb_4
XANTENNA__06639__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07485_ top.a1.instruction\[26\] net528 _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10159__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1076_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09948__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ _04276_ _04277_ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__o21ai_1
X_06436_ _01476_ _01561_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06367_ net905 net904 top.a1.instruction\[6\] _01474_ vssd1 vssd1 vccd1 vccd1 _01494_
+ sky130_fd_sc_hd__and4b_2
X_09155_ top.pc\[5\] _02641_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08106_ _03229_ _03232_ net278 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06298_ net1106 net824 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__and2_4
XFILLER_0_4_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09086_ _01584_ _01606_ _02187_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08037_ _03157_ _03163_ _01570_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06811__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold840 top.DUT.register\[15\]\[19\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 top.DUT.register\[16\]\[11\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 top.DUT.register\[10\]\[15\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 top.ramaddr\[8\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 top.DUT.register\[25\]\[17\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 top.DUT.register\[10\]\[25\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ net1699 net164 net431 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__mux2_1
X_08939_ top.pad.button_control.r_counter\[5\] top.pad.button_control.r_counter\[6\]
+ top.pad.button_control.r_counter\[7\] vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11950_ _05817_ _05819_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_106_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07524__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net2192 net141 net347 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XANTENNA__06878__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ net129 _05749_ top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ clknet_leaf_75_clk net1162 net1088 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
X_10832_ net2181 net159 net356 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08328__A _02685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07232__A _02339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13551_ clknet_leaf_71_clk _01115_ net1095 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10069__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ net171 net1755 net374 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ clknet_leaf_61_clk _00069_ net1101 vssd1 vssd1 vccd1 vccd1 top.ramstore\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13482_ clknet_leaf_38_clk _01046_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ net204 net2247 net379 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12433_ clknet_leaf_92_clk top.ru.next_FetchedData\[17\] net1000 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_191_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09044__A3 _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07055__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12364_ top.pad.button_control.r_counter\[14\] top.pad.button_control.r_counter\[13\]
+ _06144_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11315_ top.a1.dataIn\[25\] top.a1.dataIn\[24\] vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nand2_1
X_12295_ _01445_ _06071_ _06104_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__and3_1
X_11246_ top.a1.row1\[8\] _05108_ _05120_ top.a1.row2\[40\] _05125_ vssd1 vssd1 vccd1
+ vccd1 _05126_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10532__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ top.a1.dataInTemp\[10\] top.a1.data\[10\] net799 vssd1 vssd1 vccd1 vccd1
+ _05076_ sky130_fd_sc_hd__mux2_1
X_10128_ net1683 net146 net462 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13084__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12792__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ net156 net2159 net424 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__mux2_1
XANTENNA__11311__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13818_ clknet_leaf_63_clk _01359_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13749_ clknet_leaf_91_clk _01292_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[34\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07270_ top.DUT.register\[28\]\[14\] net653 net605 top.DUT.register\[18\]\[14\] _02383_
+ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a221o_1
XANTENNA__08491__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07294__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06221_ _01432_ _01434_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13298__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10707__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06152_ top.lcd.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07046__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 top.pad.button_control.noisy vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11111__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold114 top.ramstore\[4\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _01188_ vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold136 top.DUT.register\[16\]\[24\] vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 top.ramstore\[1\] vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold158 top.DUT.register\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _04891_ _04894_ _04902_ _01586_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a31o_1
Xhold169 top.ramstore\[29\] vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout605 _01668_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_8
Xfanout616 _01664_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout627 net630 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10442__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _03898_ net343 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__nand2_1
Xfanout638 _01652_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout649 _01642_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_4
X_09773_ _04769_ _04772_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__or3_1
X_06985_ top.DUT.register\[28\]\[20\] net653 net783 top.DUT.register\[31\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout284_A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _03331_ _03819_ _03830_ _03334_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_198_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08655_ _03722_ _03764_ net280 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout451_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ net283 _02731_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__nor2_1
X_08586_ _03693_ _03698_ net519 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07537_ top.DUT.register\[20\]\[4\] net749 net733 top.DUT.register\[19\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ top.DUT.register\[20\]\[5\] net747 net720 top.DUT.register\[14\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
XANTENNA__07285__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ net500 _02471_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__or2_1
X_06419_ top.DUT.register\[1\]\[30\] net686 net681 top.DUT.register\[7\]\[30\] _01545_
+ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a221o_1
XANTENNA__10617__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ top.DUT.register\[29\]\[7\] net664 net620 top.DUT.register\[26\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09138_ net910 top.pc\[3\] _04184_ _04198_ net897 vssd1 vssd1 vccd1 vccd1 _00084_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ _01819_ _01864_ _02782_ _03169_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__or4_1
XANTENNA__09266__X _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ net915 net1303 net853 _05036_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12080_ _05911_ _05946_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__nor2_2
XANTENNA__08611__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 top.DUT.register\[25\]\[27\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13524__RESET_B net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 top.DUT.register\[31\]\[22\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 top.DUT.register\[15\]\[2\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net10 net831 net830 net1333 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__a22o_1
XANTENNA__09426__B top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ clknet_leaf_2_clk _00546_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07514__X _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _05776_ _05781_ _05786_ _05790_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09161__B _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ top.a1.dataIn\[5\] _05729_ _05731_ _05732_ _05693_ vssd1 vssd1 vccd1 vccd1
+ _05734_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_129_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13603_ clknet_leaf_95_clk _01162_ net990 vssd1 vssd1 vccd1 vccd1 top.ramload\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ top.DUT.register\[28\]\[11\] net221 net356 vssd1 vssd1 vccd1 vccd1 _00997_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ _05610_ _05635_ _05638_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_31_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ clknet_leaf_15_clk _01098_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10746_ net241 net1943 net373 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__B1 _04689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13465_ clknet_leaf_36_clk _01029_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10527__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10677_ net260 net2216 net377 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07028__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08225__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ clknet_leaf_96_clk top.ru.next_FetchedData\[0\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13396_ clknet_leaf_45_clk _00960_ net1099 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09422__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__A2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ _01403_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07984__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ top.lcd.cnt_20ms\[15\] top.lcd.cnt_20ms\[14\] _06091_ top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__a31o_1
XANTENNA__10262__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11229_ net879 net880 _05098_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07736__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07200__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11882__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ top.DUT.register\[4\]\[25\] net566 net554 top.DUT.register\[7\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire517_A _01885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ net311 _03204_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08371_ _02589_ _02889_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07322_ net503 _02447_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07267__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07253_ _02363_ _02365_ _02371_ _02379_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__or4_4
XANTENNA__10437__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06204_ top.busy_o top.ru.state\[4\] vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07019__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07184_ top.DUT.register\[11\]\[13\] net642 net629 top.DUT.register\[9\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06778__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08519__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _04939_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_4
XANTENNA__09716__A1 _03616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 _04931_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_6
XANTENNA__10172__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout424 _04925_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08150__B _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_8
Xfanout446 _04950_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_4
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _04823_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__or2_1
Xfanout468 _03339_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout666_A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 _03255_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _03733_ net342 _04759_ _04763_ net339 vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__o221a_1
XANTENNA__10900__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ top.DUT.register\[27\]\[20\] net778 net725 top.DUT.register\[17\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
X_08707_ net1332 net837 net816 _03814_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__a22o_1
X_09687_ top.a1.dataIn\[5\] net794 net803 top.pc\[5\] _04704_ vssd1 vssd1 vccd1 vccd1
+ _04705_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ top.DUT.register\[20\]\[22\] net579 net645 top.DUT.register\[17\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _03648_ _03748_ net304 vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08569_ net310 _03478_ _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o21ai_4
XANTENNA_clkbuf_4_0__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ net187 net2032 net387 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07258__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11580_ _05436_ _05447_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10531_ net1983 net218 net361 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10347__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ clknet_leaf_49_clk _00814_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ net197 net1434 net371 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12201_ _05961_ _04976_ net847 top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 _01286_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_122_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ clknet_leaf_105_clk _00745_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10393_ net219 net1604 net329 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__mux2_1
X_12132_ _05994_ _05998_ _06000_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07430__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06413__X _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10082__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ _05896_ _05909_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__or3_1
XANTENNA__09156__B _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net2 net842 net812 net1340 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__o22a_1
Xfanout980 net39 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10810__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout991 net996 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ clknet_leaf_120_clk _00529_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11916_ net129 _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_142_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07497__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12896_ clknet_leaf_49_clk _00460_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09891__B1 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11847_ _05715_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ _05621_ _05638_ _05625_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09111__S _04145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ clknet_leaf_32_clk _01081_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ net185 net1760 net383 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XANTENNA__10257__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13448_ clknet_leaf_34_clk _01012_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload12 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_42_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload23 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload23/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__06209__B1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload34 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload34/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload45 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08749__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload56 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_2
X_13379_ clknet_leaf_50_clk _00943_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload67 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__clkinv_2
Xclkload78 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08522__Y _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07957__B1 _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload89 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_wire467_A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07421__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08251__A _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_11__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ top.DUT.register\[17\]\[16\] net644 net544 top.DUT.register\[5\]\[16\] _03066_
+ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07709__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ top.DUT.register\[6\]\[17\] net763 net735 top.DUT.register\[24\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_79_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09610_ _01604_ _04632_ _04639_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ net808 _01948_ net463 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__o21a_1
XANTENNA__10720__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ net529 _04576_ _04423_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__o21ai_2
X_06753_ top.DUT.register\[14\]\[25\] net721 net668 top.DUT.register\[5\]\[25\] _01879_
+ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a221o_1
XANTENNA__11117__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _04495_ _04509_ _04510_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__and3_1
XANTENNA__07488__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06684_ top.DUT.register\[25\]\[27\] net623 net540 top.DUT.register\[22\]\[27\] _01810_
+ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a221o_1
XANTENNA__09882__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ net314 net490 vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nand2_2
XANTENNA__06696__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__D net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08354_ _03314_ _03323_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07305_ top.DUT.register\[11\]\[9\] net640 net557 top.DUT.register\[6\]\[9\] _02431_
+ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ net298 _03127_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__nand2_2
Xclkload6 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__10167__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout414_A _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09956__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07236_ top.DUT.register\[26\]\[14\] net761 net691 top.DUT.register\[3\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ top.DUT.register\[1\]\[13\] net687 _02288_ _02293_ vssd1 vssd1 vccd1 vccd1
+ _02294_ sky130_fd_sc_hd__a211o_1
X_07098_ _02216_ _02218_ _02220_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06620__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__A2_N _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 _04738_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout221 _04732_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 _04726_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout243 _04711_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08960__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout254 _04703_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
X_09808_ _03832_ net340 net337 _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__o211a_4
XANTENNA__10630__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout298 net301 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ net199 net1772 net439 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12750_ clknet_leaf_110_clk _00314_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08676__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07479__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11701_ _05568_ _05569_ _05565_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__a21o_1
XFILLER_0_194_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06687__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12681_ clknet_leaf_3_clk _00245_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11632_ _05409_ _05471_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__nor2_1
XANTENNA__08428__A1 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06408__X _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11563_ _05430_ _05432_ _05395_ _05428_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10077__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08055__B _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ clknet_leaf_120_clk _00866_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10514_ net1944 net151 net361 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__mux2_1
X_11494_ _05338_ _05352_ _05362_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09389__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ clknet_leaf_12_clk _00797_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10445_ net145 net2249 net324 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
XANTENNA__10805__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07403__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13164_ clknet_leaf_8_clk _00728_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08071__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ net445 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__inv_2
XANTENNA__08600__B2 _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06611__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _05977_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__or2_1
X_13095_ clknet_leaf_8_clk _00659_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12046_ _05902_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08364__B1 _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09313__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ clknet_leaf_62_clk _00512_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08667__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__B2 _03776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12879_ clknet_leaf_22_clk _00443_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08419__B2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07890__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08246__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08070_ _03193_ _03196_ net276 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload101 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_12
XANTENNA__07642__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07021_ top.DUT.register\[13\]\[11\] net649 net606 top.DUT.register\[18\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
XANTENNA__06850__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10715__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09077__A _01909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ _02033_ net592 net1222 net868 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09805__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ top.DUT.register\[27\]\[16\] net776 net678 top.DUT.register\[13\]\[16\] _03049_
+ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__a221o_1
Xhold18 _01182_ vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 _01191_ vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__Y _04145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ top.DUT.register\[20\]\[18\] net579 net666 top.DUT.register\[29\]\[18\] _02980_
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10450__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ top.DUT.register\[14\]\[24\] net614 net596 top.DUT.register\[27\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07785_ top.DUT.register\[20\]\[19\] net749 net714 top.DUT.register\[30\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a22o_1
XANTENNA__08107__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_A _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ _04559_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_84_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08658__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06736_ _01840_ _01859_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_203_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07612__X _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ _04494_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__nand2_1
XANTENNA__12377__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ top.DUT.register\[15\]\[27\] net704 _01791_ _01793_ vssd1 vssd1 vccd1 vccd1
+ _01794_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout629_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08406_ _02891_ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__xnor2_1
X_09386_ _04422_ _04429_ _01619_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__a21o_1
XANTENNA__08156__A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07881__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06598_ top.DUT.register\[14\]\[29\] net614 _01715_ _01722_ _01724_ vssd1 vssd1 vccd1
+ vccd1 _01725_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_62_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08337_ net476 _03452_ _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07094__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08830__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ net1376 net837 net816 _03392_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a22o_1
XANTENNA__07633__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout998_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06841__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07219_ top.DUT.register\[7\]\[15\] net552 net624 top.DUT.register\[25\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10625__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ _03323_ _03324_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_197_Right_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10230_ net154 net2094 net407 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ net157 net1738 net415 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1005 net1008 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1019 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_2
Xfanout1027 net1029 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_4
X_10092_ net160 net2128 net417 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
Xfanout1038 net1051 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10360__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13851_ net1116 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_199_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ clknet_leaf_42_clk _00366_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13782_ clknet_leaf_64_clk _01325_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10994_ net1436 _05011_ net535 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12733_ clknet_leaf_108_clk _00297_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12664_ clknet_leaf_107_clk _00228_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07872__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ _05482_ _05483_ top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11204__B _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ clknet_leaf_5_clk _00159_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12749__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ _05413_ _05415_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nor2_1
XANTENNA__07624__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06832__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10535__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ _05341_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire496 _02779_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
X_13216_ clknet_leaf_42_clk _00780_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ net200 net1693 net326 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__mux2_1
XANTENNA__09377__A2 _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ clknet_leaf_52_clk _00711_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10359_ net1530 net186 net394 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ clknet_leaf_121_clk _00642_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_183_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _05897_ _05898_ _05885_ _05895_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a211o_1
XANTENNA__10270__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06899__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ top.DUT.register\[6\]\[3\] net556 net544 top.DUT.register\[5\]\[3\] _02693_
+ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ _01590_ _01631_ _01643_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_66_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09240_ top.pc\[11\] _04280_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__and2_1
X_06452_ top.a1.instruction\[13\] net820 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__or2_1
XANTENNA__07863__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09171_ top.pc\[6\] _02612_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nand2b_1
X_06383_ top.a1.instruction\[19\] _01498_ _01499_ vssd1 vssd1 vccd1 vccd1 _01510_
+ sky130_fd_sc_hd__and3_4
XFILLER_0_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06990__Y _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06208__B top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08122_ net499 net294 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__nand2_1
XANTENNA__09736__A1_N net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07615__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08053_ _03165_ _03172_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__nand2_1
XANTENNA__10445__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__B net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ top.DUT.register\[2\]\[11\] net717 _02129_ _02130_ vssd1 vssd1 vccd1 vccd1
+ _02131_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08576__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ net497 net591 net1351 net865 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06511__X _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout579_A _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _03012_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and2_1
XANTENNA__10180__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08886_ net270 _03841_ _03982_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07000__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ top.DUT.register\[7\]\[18\] net682 _02958_ _02963_ vssd1 vssd1 vccd1 vccd1
+ _02964_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout746_A _01518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A1_N _03183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ net499 _02492_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__and2b_1
XFILLER_0_195_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _04519_ _04522_ _04520_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a21bo_1
X_06719_ top.DUT.register\[2\]\[26\] net661 net570 top.DUT.register\[8\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07699_ top.DUT.register\[10\]\[0\] net727 net674 top.DUT.register\[18\]\[0\] _02825_
+ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_121_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08500__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09438_ _04477_ _04478_ _01618_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07854__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09369_ top.pc\[18\] _04385_ top.pc\[19\] vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _05232_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12380_ clknet_leaf_70_clk top.edg2.button_i net1105 vssd1 vssd1 vccd1 vccd1 top.edg2.flip1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _05185_ _05192_ _05194_ _05200_ top.a1.dataIn\[25\] vssd1 vssd1 vccd1 vccd1
+ _05201_ sky130_fd_sc_hd__o32a_1
XANTENNA__06814__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11262_ top.a1.row1\[2\] _05094_ _05107_ top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1
+ _05140_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13001_ clknet_leaf_3_clk _00565_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10213_ net209 net2162 net407 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__mux2_1
X_11193_ net850 _05070_ net531 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__and3_1
X_10144_ net220 net1811 net415 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08319__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06593__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10090__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ net224 net1564 net418 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ clknet_leaf_68_clk _01375_ net1106 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13765_ clknet_leaf_74_clk _01308_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10977_ top.a1.halfData\[2\] net797 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11215__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12716_ clknet_leaf_9_clk _00280_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07845__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13696_ clknet_leaf_75_clk _01244_ net1088 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09047__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ clknet_leaf_7_clk _00211_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12578_ clknet_leaf_43_clk _00142_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06805__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11529_ _05381_ _05387_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10265__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 top.DUT.register\[14\]\[27\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 top.DUT.register\[11\]\[18\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold329 top.DUT.register\[11\]\[14\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08530__Y _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 _01562_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_4
XANTENNA__09123__A_N net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06584__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1007 top.DUT.register\[10\]\[7\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07146__Y _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ _02080_ _03090_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__xnor2_2
Xhold1018 top.DUT.register\[15\]\[22\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 top.DUT.register\[29\]\[23\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11226__A_N net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08671_ _02993_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07622_ top.DUT.register\[9\]\[2\] net627 net607 top.DUT.register\[12\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07553_ top.DUT.register\[15\]\[4\] net706 net680 top.DUT.register\[13\]\[4\] _02679_
+ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06504_ net900 net801 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nand2_2
XANTENNA__11125__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07322__B _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ _02563_ _02609_ _02206_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_200_Right_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ net137 _04269_ _04274_ net819 net909 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__o221a_1
X_06435_ _01476_ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout327_A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07049__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ _04200_ _04203_ _04202_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__a21o_1
X_06366_ _01426_ _01427_ net866 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_79_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08105_ _03230_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10175__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ _01609_ _03153_ _04146_ _01489_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__o2bb2a_1
X_06297_ net1104 _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__and2_4
XFILLER_0_140_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09964__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ net903 net901 top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or3b_1
XANTENNA__09817__X _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold830 top.DUT.register\[5\]\[26\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold841 top.DUT.register\[6\]\[13\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold852 wb.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12524__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 top.DUT.register\[10\]\[5\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10903__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 top.DUT.register\[17\]\[19\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 top.DUT.register\[31\]\[4\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 top.DUT.register\[19\]\[27\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07221__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ net1961 net168 net430 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout863_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06575__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ top.pad.button_control.r_counter\[10\] top.pad.button_control.r_counter\[9\]
+ top.pad.button_control.r_counter\[7\] top.pad.button_control.r_counter\[5\] vssd1
+ vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nand4_1
XANTENNA__09552__X _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ _03237_ _03825_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net1732 net146 net346 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11880_ net129 _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10831_ net1536 net160 net353 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08328__B _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ clknet_leaf_69_clk _01114_ net1104 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07288__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10762_ net178 net2007 net373 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__mux2_1
XANTENNA__07827__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ clknet_leaf_114_clk _00068_ net939 vssd1 vssd1 vccd1 vccd1 top.ramstore\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13481_ clknet_leaf_4_clk _01045_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10693_ net214 net1314 net379 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08615__Y _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ clknet_leaf_92_clk top.ru.next_FetchedData\[16\] net1000 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[16\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_33_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06416__X _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10085__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12363_ _06146_ _06147_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11314_ top.a1.dataIn\[31\] top.a1.dataIn\[30\] _05183_ vssd1 vssd1 vccd1 vccd1 _05184_
+ sky130_fd_sc_hd__nand3_1
XANTENNA__09727__X _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ top.lcd.cnt_500hz\[5\] _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08631__X _03742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09737__C1 _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ net891 top.a1.row1\[112\] _05105_ _05100_ _01444_ vssd1 vssd1 vccd1 vccd1
+ _05125_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10813__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09175__A _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11176_ net1288 net532 net525 _05075_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a22o_1
X_10127_ net1551 net155 net460 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ net161 net2278 net421 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13817_ clknet_leaf_70_clk _01358_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap494_A _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13053__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07279__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13748_ clknet_leaf_88_clk _01291_ net1005 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[33\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07818__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13679_ clknet_leaf_94_clk _00006_ net993 vssd1 vssd1 vccd1 vccd1 top.ru.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06220_ _01434_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
XANTENNA__08254__A _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09440__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 net84 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07451__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold115 _01171_ vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 top.a1.row1\[60\] vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold137 top.a1.dataInTemp\[8\] vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 top.DUT.register\[9\]\[7\] vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09910_ _04891_ _04894_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a21oi_1
Xhold159 top.DUT.register\[28\]\[14\] vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10723__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 _01668_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_4
X_09841_ net175 top.DUT.register\[1\]\[23\] net437 vssd1 vssd1 vccd1 vccd1 _00145_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07203__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout617 _01664_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_60_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout628 net630 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 _01648_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_4
XANTENNA__06557__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__B1 _02854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _04776_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nor2_1
X_06984_ top.DUT.register\[21\]\[20\] net574 net601 top.DUT.register\[10\]\[20\] _02110_
+ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a221o_1
X_08723_ _02121_ _03086_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_198_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08703__B1 _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ _03275_ _03299_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nand2_1
XANTENNA__07604__Y _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08429__A _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ net283 _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__and2_1
X_08585_ _03496_ _03541_ _03585_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10030__Y _04925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09259__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout444_A _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ net806 _02641_ _02661_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__o21a_1
XANTENNA__09959__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07467_ top.DUT.register\[17\]\[5\] _01520_ net735 top.DUT.register\[24\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout611_A _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ _02516_ _02521_ _04250_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__o21ba_1
X_06418_ top.DUT.register\[8\]\[30\] net739 net711 top.DUT.register\[9\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a22o_1
XANTENNA__08164__A _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ top.DUT.register\[25\]\[7\] net623 net540 top.DUT.register\[22\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09137_ net133 _04191_ _04197_ net910 vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_134_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06349_ net903 net902 net901 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__a21o_2
XFILLER_0_71_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07442__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ _03414_ _04124_ _04126_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout980_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06796__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ _03141_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__nor2_4
XANTENNA__10633__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 top.DUT.register\[30\]\[2\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 top.DUT.register\[15\]\[8\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold682 top.DUT.register\[26\]\[17\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net9 net841 net811 net1280 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__o22a_1
XANTENNA__07508__A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 top.DUT.register\[21\]\[31\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06548__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ clknet_leaf_4_clk _00545_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11932_ _05797_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11863_ _05731_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06720__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13602_ clknet_leaf_95_clk _01161_ net990 vssd1 vssd1 vccd1 vccd1 top.ramload\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10814_ net1400 net223 net353 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _05635_ _05638_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10745_ net244 net1973 net376 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__mux2_1
X_13533_ clknet_leaf_107_clk _01097_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09670__A1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10808__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__B2 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06484__A1 top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ clknet_leaf_111_clk _01028_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08074__A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10676_ net263 net1584 net379 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ clknet_leaf_94_clk top.ru.next_dready net992 vssd1 vssd1 vccd1 vccd1 top.d_ready
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08225__A2 _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ clknet_leaf_5_clk _00959_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12346_ net2222 _06134_ _06136_ net796 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__o211a_1
XANTENNA__07433__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06787__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ net1248 _06092_ _06094_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10543__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__S _04145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11228_ net882 net884 _05093_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_1
XFILLER_0_208_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ net1349 net532 _05065_ _05067_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__a22o_1
XANTENNA_max_cap507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06711__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ net1304 net838 net817 _03491_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a22o_1
XANTENNA__06992__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ net503 _02447_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__and2_1
XFILLER_0_190_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10718__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ _02373_ _02375_ _02376_ _02378_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__or4_1
XANTENNA__07672__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06203_ _00008_ top.a1.nextHex\[7\] vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[4\] sky130_fd_sc_hd__or2_1
X_07183_ top.DUT.register\[5\]\[13\] net546 net543 top.DUT.register\[22\]\[13\] _02309_
+ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07424__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06778__A2 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07975__A1 _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10453__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09716__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 _04939_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_8
Xfanout414 _04931_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_4
Xfanout425 net428 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_8
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _04918_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09824_ _04813_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__nor2_1
Xfanout447 net449 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1101_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout469 _03339_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
XANTENNA__09543__A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06967_ top.DUT.register\[30\]\[20\] net714 net677 top.DUT.register\[18\]\[20\] _02091_
+ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a221o_1
X_09755_ _01586_ _04761_ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout561_A _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09262__B _04304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net888 top.pc\[19\] net538 _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__a22o_1
XANTENNA__11287__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ net836 _04212_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08159__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06898_ top.DUT.register\[26\]\[22\] net622 net613 top.DUT.register\[14\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09830__X _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08637_ net278 _03700_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_194_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ net285 _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__or2_1
XANTENNA__12957__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08446__X _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07519_ top.DUT.register\[13\]\[4\] net650 net645 top.DUT.register\[17\]\[4\] _02645_
+ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08499_ _03601_ _03609_ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nand3_2
XANTENNA__10628__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ net1658 net227 net362 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07663__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10461_ net201 top.DUT.register\[17\]\[13\] net372 vssd1 vssd1 vccd1 vccd1 _00647_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12200_ net2345 net845 net813 _05975_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ clknet_leaf_56_clk _00744_ net1086 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10392_ net224 net2283 net327 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__mux2_1
XANTENNA__06769__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__A1 _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ _05994_ _05998_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__o21a_1
XANTENNA__10363__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12062_ _05920_ _05921_ _05918_ _05919_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a211o_1
XANTENNA__09707__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 top.DUT.register\[14\]\[26\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ top.busy_o net831 wb.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__or3b_1
XANTENNA__08391__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net979 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07194__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09453__A _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout992 net995 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06941__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12964_ clknet_leaf_39_clk _00528_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1190 top.DUT.register\[21\]\[0\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_11915_ _05745_ _05753_ _05743_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a21o_1
XANTENNA__06205__B1_N top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ clknet_leaf_113_clk _00459_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11846_ _05689_ net130 _05679_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _05621_ _05625_ _05638_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__and3_1
XANTENNA__10538__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13516_ clknet_leaf_10_clk _01080_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10728_ net188 net2080 net383 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10659_ net1736 net227 net453 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
X_13447_ clknet_leaf_8_clk _01011_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_8
Xclkload24 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__06209__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload35 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload35/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload46 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__07406__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ clknet_leaf_43_clk _00942_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08532__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload57 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_12
XANTENNA__06604__X _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload68 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_2
Xclkload79 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinv_4
X_12329_ top.pad.button_control.r_counter\[0\] net1231 _06125_ vssd1 vssd1 vccd1 vccd1
+ _01354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10273__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07148__A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__X _04908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07870_ top.DUT.register\[29\]\[17\] net700 net696 top.DUT.register\[23\]\[17\] _02996_
+ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08382__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07185__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ _01943_ _01945_ _01946_ _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__nor4_2
XANTENNA__06932__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09540_ top.a1.instruction\[28\] net822 _04540_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__o21a_1
X_06752_ top.DUT.register\[24\]\[25\] net736 net705 top.DUT.register\[15\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ _04495_ _04510_ _04509_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06683_ top.DUT.register\[1\]\[27\] net655 net552 top.DUT.register\[7\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ net317 net310 vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__nand2_4
XANTENNA__07893__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__X _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07170__X _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08353_ net314 _03470_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10448__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout142_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07304_ top.DUT.register\[29\]\[9\] net664 net624 top.DUT.register\[25\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_178_Right_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08284_ _03284_ _03291_ net286 vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__mux2_1
XANTENNA__07645__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_46_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06999__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07235_ top.DUT.register\[28\]\[14\] net586 net687 top.DUT.register\[1\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10972__A top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07166_ top.DUT.register\[7\]\[13\] net682 net672 top.DUT.register\[16\]\[13\] _02292_
+ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a221o_1
XANTENNA__09538__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10183__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07097_ top.DUT.register\[2\]\[10\] net660 net604 top.DUT.register\[18\]\[10\] _02223_
+ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__A top.a1.instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09972__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net202 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout776_A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 _04732_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_1
Xfanout233 _04726_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13430__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10911__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 net258 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07176__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _04693_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
X_09807_ net802 _04807_ _04808_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a211o_1
Xfanout288 _02855_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
Xfanout299 net301 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ _03110_ _03111_ _03117_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nor4_1
XFILLER_0_199_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09738_ _03689_ net341 net338 _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_2_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09669_ net149 net2196 net437 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11700_ _05568_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__nand2_1
X_12680_ clknet_leaf_33_clk _00244_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12209__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ _05470_ _05471_ _05482_ _05483_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a22o_1
XANTENNA__10358__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11562_ _05426_ _05431_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07100__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ net465 _04919_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__nor2_4
X_13301_ clknet_leaf_7_clk _00865_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _05353_ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13232_ clknet_leaf_0_clk _00796_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ net155 net1585 net325 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10093__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ clknet_leaf_29_clk _00727_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10375_ _01601_ net465 _04929_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__nor3_4
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12114_ _05974_ _05975_ _05979_ _05983_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__o22a_2
X_13094_ clknet_leaf_14_clk _00658_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ _05887_ _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nor2_1
XANTENNA__10821__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08364__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__B2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06914__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_2_clk _00511_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12878_ clknet_leaf_117_clk _00442_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11829_ _05659_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload102 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__clkinvlp_4
X_07020_ top.DUT.register\[2\]\[11\] net661 net543 top.DUT.register\[22\]\[11\] _02146_
+ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09077__B _02879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12215__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08971_ _02075_ net591 net1346 net868 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__a2bb2o_1
X_07922_ top.DUT.register\[26\]\[16\] net760 net716 top.DUT.register\[2\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a22o_1
XANTENNA__10731__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 top.a1.dataInTemp\[5\] vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__A _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ top.DUT.register\[21\]\[18\] net574 net606 top.DUT.register\[18\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__a22o_1
XANTENNA__07606__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__A1_N net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06905__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ top.DUT.register\[3\]\[24\] net788 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__and2_1
X_07784_ top.DUT.register\[19\]\[19\] net734 _01535_ top.DUT.register\[3\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09380__X _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__A top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09523_ _01840_ _04542_ _04546_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_84_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06735_ _01840_ _01859_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_203_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10967__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout357_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _01991_ _04493_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06666_ top.DUT.register\[30\]\[27\] net712 net681 top.DUT.register\[7\]\[27\] _01792_
+ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a221o_1
XANTENNA__06509__X _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07330__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08405_ _03523_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__nand2_2
XFILLER_0_148_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10178__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09385_ _04422_ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06597_ top.DUT.register\[11\]\[29\] net641 net542 top.DUT.register\[22\]\[29\] _01723_
+ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_191_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08336_ net482 net275 _03456_ _03453_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__o31a_1
XANTENNA__07618__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09967__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08267_ net887 net895 net536 _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a22o_1
XANTENNA__10906__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ top.DUT.register\[9\]\[15\] net627 net548 top.DUT.register\[24\]\[15\] _02344_
+ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08172__A _02339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ _02562_ net289 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07149_ net508 _02274_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_95_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11310__B net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07397__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ net161 net2284 net414 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1008 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
X_10091_ net164 net1968 net420 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10641__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 net1019 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
Xfanout1039 net1042 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13850_ net1115 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12801_ clknet_leaf_23_clk _00365_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13781_ clknet_leaf_64_clk _01324_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10993_ top.a1.dataIn\[6\] net848 net843 _05010_ vssd1 vssd1 vccd1 vccd1 _05011_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07857__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ clknet_leaf_18_clk _00296_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13326__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10088__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ clknet_leaf_77_clk _00227_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _05482_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ clknet_leaf_48_clk _00158_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11545_ _05380_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10816__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__Y _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11476_ _05325_ _05332_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08082__A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ clknet_leaf_113_clk _00779_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10427_ net209 net2264 net325 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10916__A0 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10358_ net1942 net187 net394 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ clknet_leaf_15_clk _00710_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06596__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10551__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ clknet_leaf_10_clk _00641_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10289_ net1713 net194 net404 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__mux2_1
XANTENNA__08337__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _05874_ _05876_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_183_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2__f_clk_X clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06520_ _01573_ net789 _01634_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_66_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07848__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07312__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06451_ _01388_ net820 _01576_ _01571_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09170_ _04213_ _04216_ _04215_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06382_ _01499_ net791 _01506_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__and3_4
X_08121_ _03246_ _03247_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10726__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ _03165_ _03172_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07003_ top.DUT.register\[31\]\[11\] net746 net715 top.DUT.register\[30\]\[11\] _02128_
+ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08974__A2_N net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07379__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08576__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08576__B2 _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06587__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10461__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09535__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ net1274 net870 _02660_ net593 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__a22o_1
XANTENNA__08359__A2_N _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ net807 _03031_ _01624_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_205_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08885_ net300 _03904_ net274 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout474_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ top.DUT.register\[18\]\[18\] net677 net670 top.DUT.register\[5\]\[18\] _02962_
+ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13349__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__inv_2
XFILLER_0_196_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout739_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__Y _02469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _01840_ _04542_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__xor2_1
XANTENNA__07839__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06718_ top.DUT.register\[11\]\[26\] net641 net546 top.DUT.register\[5\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
X_07698_ top.DUT.register\[25\]\[0\] net771 net763 top.DUT.register\[6\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07303__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08500__B2 _03616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _04477_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06649_ _01755_ _01774_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ top.pc\[18\] top.pc\[19\] _04385_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13518__RESET_B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07067__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ net268 _03440_ _03441_ net272 _03439_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_97_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_113_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09299_ _01615_ _02688_ _02736_ net823 _01622_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__o221a_4
XANTENNA__10636__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10071__A0 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13__f_clk_X clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _05189_ _05193_ _05192_ _01392_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_151_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ net891 top.a1.row1\[114\] _05105_ _05138_ vssd1 vssd1 vccd1 vccd1 _05139_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08016__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10212_ net220 net2200 net407 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__mux2_1
X_13000_ clknet_leaf_35_clk _00564_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11192_ net850 _05069_ net531 _05083_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a31o_1
XANTENNA__08630__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ net225 net1629 net414 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XANTENNA__08319__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ net232 net1419 net418 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
XANTENNA__07542__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__X _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ clknet_leaf_68_clk _01374_ net1106 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06750__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13764_ clknet_leaf_85_clk _01307_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10976_ top.a1.data\[1\] _04998_ _04989_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11215__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12715_ clknet_leaf_30_clk _00279_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13695_ clknet_leaf_71_clk _01243_ net1095 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[111\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_139_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12646_ clknet_leaf_24_clk _00210_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09047__A2 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12577_ clknet_leaf_28_clk _00141_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11528_ _05368_ _05394_ _05395_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__and4b_1
XFILLER_0_159_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 top.DUT.register\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08007__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold319 top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
X_11459_ _05326_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_185_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07708__X _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06569__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13129_ clknet_leaf_4_clk _00693_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10281__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__C_N top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__X _04915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 top.DUT.register\[1\]\[27\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 top.DUT.register\[29\]\[12\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08670_ _03737_ _03778_ _03033_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08539__X _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08730__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09371__A top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07621_ top.DUT.register\[1\]\[2\] net655 net564 top.DUT.register\[4\]\[2\] _02747_
+ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06741__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ top.DUT.register\[30\]\[4\] net714 net702 top.DUT.register\[29\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06503_ net900 net801 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07483_ top.a1.instruction\[17\] _01617_ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07297__B2 top.a1.instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11125__B net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06434_ net905 net904 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__nand2_1
X_09222_ _04258_ _04260_ _04275_ net134 vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09153_ _04210_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nand2b_1
X_06365_ top.d_ready _01489_ _01490_ top.ru.next_read_i vssd1 vssd1 vccd1 vccd1 _00007_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout222_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06506__Y _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ _02608_ net289 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _01584_ _01606_ net903 vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a21oi_1
X_06296_ net824 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
X_08035_ net490 _03148_ _03154_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__o211a_1
XANTENNA__13021__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 top.DUT.register\[6\]\[5\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 top.DUT.register\[16\]\[4\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 top.DUT.register\[16\]\[16\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold853 top.DUT.register\[26\]\[11\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold864 top.DUT.register\[10\]\[31\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 top.DUT.register\[17\]\[2\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 top.DUT.register\[12\]\[19\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 top.DUT.register\[16\]\[5\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ net1380 net171 net432 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09980__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ top.pad.button_control.r_counter\[14\] top.pad.button_control.r_counter\[13\]
+ top.pad.button_control.r_counter\[12\] top.pad.button_control.r_counter\[11\] vssd1
+ vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__or4_1
XANTENNA__06980__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ net322 _03651_ _03966_ net274 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__o22ai_1
XANTENNA__08721__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07819_ _02931_ _02933_ _02945_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__or3_1
XFILLER_0_211_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ _01909_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06732__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ net1828 net165 net356 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09277__A2 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10761_ net183 net1781 net376 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ clknet_leaf_75_clk _00067_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13480_ clknet_leaf_34_clk _01044_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10692_ net215 net2340 net377 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12431_ clknet_leaf_93_clk top.ru.next_FetchedData\[15\] net999 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10366__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08788__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ net2090 _06144_ net795 vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08912__X _04009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06799__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11313_ top.a1.dataIn\[27\] top.a1.dataIn\[26\] top.a1.dataIn\[29\] top.a1.dataIn\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or4_1
X_12293_ _06098_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11244_ top.a1.row1\[56\] _05112_ _05116_ top.a1.row1\[104\] _05123_ vssd1 vssd1
+ vccd1 vccd1 _05124_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09175__B _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ top.a1.dataInTemp\[9\] top.a1.data\[9\] net799 vssd1 vssd1 vccd1 vccd1 _05075_
+ sky130_fd_sc_hd__mux2_1
X_10126_ net1311 net158 net460 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08960__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10057_ net164 net1990 net424 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11311__A3 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06723__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ clknet_leaf_70_clk _01357_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13747_ clknet_leaf_87_clk _01290_ net1008 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[32\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08476__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959_ net1290 _04979_ _04986_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13678_ clknet_leaf_94_clk _00011_ net993 vssd1 vssd1 vccd1 vccd1 top.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10276__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ clknet_leaf_6_clk _00193_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08228__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08254__B _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__B2 _03882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold105 _01168_ vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold116 top.ramstore\[14\] vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 top.ramload\[12\] vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 top.DUT.register\[16\]\[26\] vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07585__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold149 top.ramstore\[30\] vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 _01667_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_8
X_09840_ _03882_ net342 net339 _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__o211a_2
Xfanout618 _01664_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__buf_4
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_4
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08951__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ top.pc\[17\] _04394_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nor2_1
X_06983_ top.DUT.register\[1\]\[20\] net658 net613 top.DUT.register\[14\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a22o_1
X_08722_ net522 _03827_ _03828_ net478 vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_198_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08703__B2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ net314 _03297_ _03543_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__o21ai_2
XANTENNA__06714__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07604_ _02724_ _02730_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__nor2_8
X_08584_ _02401_ net484 net480 _03695_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ net806 _02641_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout437_A _04681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07466_ top.DUT.register\[19\]\[5\] net731 net727 top.DUT.register\[10\]\[5\] _02590_
+ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06417_ _01497_ net791 _01506_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__and3_1
X_09205_ _04257_ _04259_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08219__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ top.DUT.register\[1\]\[7\] net655 net604 top.DUT.register\[18\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout604_A _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08164__B net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06348_ net902 top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__nor2_1
X_09136_ _04159_ _04163_ _04194_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09067_ _04127_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10914__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06279_ net2352 net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[23\] sky130_fd_sc_hd__and2_1
XFILLER_0_130_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09719__B1 _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08018_ _03129_ _03142_ _03143_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__or4_1
XANTENNA__07993__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 top.DUT.register\[29\]\[6\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 top.DUT.register\[24\]\[3\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09195__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 top.DUT.register\[8\]\[25\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 top.pad.button_control.r_counter\[11\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 top.pad.button_control.r_counter\[4\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07745__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ net1722 net240 net430 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ clknet_leaf_59_clk _00544_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11931_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06705__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11046__A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ _01398_ _05684_ net130 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08907__X _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ clknet_leaf_95_clk _01160_ net988 vssd1 vssd1 vccd1 vccd1 top.ramload\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10813_ net1385 net233 net354 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11793_ _05633_ _05659_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_45_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ clknet_leaf_17_clk _01096_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10744_ net248 net1951 net373 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__mux2_1
XANTENNA__06427__X _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07130__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06484__A2 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ clknet_leaf_105_clk _01027_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10096__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ net149 net1804 net377 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12414_ clknet_leaf_94_clk net874 net997 vssd1 vssd1 vccd1 vccd1 top.i_ready sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09738__X _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13394_ clknet_leaf_48_clk _00958_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ top.pad.button_control.r_counter\[7\] _06134_ vssd1 vssd1 vccd1 vccd1 _06136_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_189_Left_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10824__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__Y _03483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07984__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ net1248 _06092_ net1107 vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11227_ net884 _05099_ net882 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_56_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07197__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07736__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output66_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ top.a1.data\[1\] net798 _04996_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06944__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ net2211 net219 net460 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
X_11089_ net66 net859 vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_198_Left_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09920__Y _04912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11048__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07320_ _02427_ net501 net807 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_2
XANTENNA__07440__Y _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ top.DUT.register\[17\]\[14\] net724 net709 top.DUT.register\[9\]\[14\] _02377_
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06202_ net1180 _01423_ _01419_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[3\] sky130_fd_sc_hd__or3b_1
XFILLER_0_54_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07182_ top.DUT.register\[29\]\[13\] net666 net618 top.DUT.register\[30\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10734__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout404 _04939_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_4
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
Xfanout426 net428 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
Xfanout437 _04681_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_8
X_09823_ _04812_ _04814_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__nor2_1
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 net462 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_6
XANTENNA_fanout387_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _04751_ _04755_ _04760_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a21oi_1
X_06966_ top.DUT.register\[14\]\[20\] net722 net682 top.DUT.register\[7\]\[20\] _02092_
+ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a221o_1
X_08705_ _03331_ _03797_ _03812_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09685_ net251 net1860 net439 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__mux2_1
X_06897_ top.DUT.register\[6\]\[22\] net559 net546 top.DUT.register\[5\]\[22\] _02023_
+ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net287 _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07360__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08567_ _03581_ _03680_ net307 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__mux2_1
XANTENNA__10909__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A _01527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_202_Left_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout819_A _01588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ top.DUT.register\[2\]\[4\] net661 net597 top.DUT.register\[27\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a22o_1
XANTENNA__08175__A _02298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07112__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ _03334_ _03596_ _03614_ net477 vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11313__B top.a1.dataIn\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07449_ top.DUT.register\[5\]\[6\] net546 net606 top.DUT.register\[18\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08860__B1 _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ net207 net1508 net369 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ _04166_ _04171_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__and2b_1
XANTENNA__07415__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ net233 net1897 net328 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10644__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _05979_ _05983_ _05996_ _05980_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07966__A2 _02034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10970__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_211_Left_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12061_ _05920_ _05921_ _05918_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 top.DUT.register\[5\]\[16\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 top.DUT.register\[17\]\[23\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07718__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ top.busy_o wb.prev_BUSY_O net842 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__and3b_1
XANTENNA__06926__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 net964 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
Xfanout971 net978 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 net986 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout993 net995 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12963_ clknet_leaf_33_clk _00527_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1180 top.DUT.register\[24\]\[17\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_84_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1191 top.pad.keyCode\[7\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11914_ _05776_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12894_ clknet_leaf_13_clk _00458_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07351__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11845_ _05679_ _05689_ net130 vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nand3_1
XANTENNA__10819__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11504__A top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11776_ _01397_ _05642_ _05643_ _05644_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13515_ clknet_leaf_30_clk _01079_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ net194 net1641 net383 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XANTENNA__08851__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ clknet_leaf_24_clk _01010_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10658_ net1404 net180 net450 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
Xclkload14 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_70_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload25 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08682__A2_N net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload36 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_6
XANTENNA__10554__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload47 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload47/X sky130_fd_sc_hd__clkbuf_8
X_13377_ clknet_leaf_28_clk _00941_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10589_ net223 net2072 net385 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
Xclkload58 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_6
XFILLER_0_152_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload69 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_140_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12328_ top.pad.button_control.r_counter\[0\] net1231 net795 vssd1 vssd1 vccd1 vccd1
+ _06125_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_167_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12259_ _06082_ _06083_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__nor2_1
XANTENNA__07148__B _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07709__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06917__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07435__Y _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ top.DUT.register\[16\]\[24\] net637 net609 top.DUT.register\[12\]\[24\] _01933_
+ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07590__B1 _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13455__RESET_B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09082__C _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06751_ top.DUT.register\[31\]\[25\] net744 net697 top.DUT.register\[23\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a22o_1
XANTENNA__11269__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_75_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09470_ _04492_ _04494_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__nand2_1
X_06682_ top.DUT.register\[5\]\[27\] net544 _01800_ _01808_ vssd1 vssd1 vccd1 vccd1
+ _01809_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_69_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08421_ net322 _02712_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__nor2_2
XFILLER_0_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06696__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08352_ net270 _03472_ _03473_ net274 vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_18_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07303_ top.DUT.register\[8\]\[9\] net571 net561 top.DUT.register\[23\]\[9\] _02429_
+ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a221o_1
XANTENNA__11133__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08283_ net285 _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload8 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07234_ _02359_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10972__B net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ top.DUT.register\[25\]\[13\] net773 net710 top.DUT.register\[9\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a22o_1
XANTENNA__10464__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06514__Y _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ top.DUT.register\[6\]\[10\] net557 net631 top.DUT.register\[19\]\[10\] _02222_
+ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_113_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06243__A top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06620__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout212 _04795_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout223 _04729_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06530__X _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout671_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _04726_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_1
Xfanout245 _04711_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout256 net258 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _04443_ net526 net332 top.a1.dataIn\[20\] net334 vssd1 vssd1 vccd1 vccd1
+ _04809_ sky130_fd_sc_hd__a221o_1
Xfanout267 _05333_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
XFILLER_0_157_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout289 net291 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_2
X_07998_ _03120_ _03122_ _03124_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__or3_1
XANTENNA__07581__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _04329_ net527 _04746_ _04718_ _04744_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__a2111o_1
X_06949_ net808 _02075_ net463 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_66_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09668_ _03261_ net342 net339 _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__o211a_2
X_08619_ _02359_ net489 _03721_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__o211a_1
XANTENNA__12209__A1 top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10639__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06687__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ _01410_ net850 _04628_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11630_ _05451_ _05494_ _05496_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__or4b_1
XFILLER_0_194_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ _05388_ net250 _05397_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__a21oi_1
X_13300_ clknet_leaf_60_clk _00864_ net1102 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10512_ net142 net1569 net367 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__mux2_1
XANTENNA__08633__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ _05358_ _05359_ _05355_ _05356_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_21_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09389__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13231_ clknet_leaf_20_clk _00795_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10443_ net158 net1700 net326 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ clknet_leaf_34_clk _00726_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ net466 _04930_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__nand2_8
X_12113_ _05967_ _05982_ _05975_ _05971_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06611__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13093_ clknet_leaf_118_clk _00657_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12044_ _05852_ _05859_ net127 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_53_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__A2 _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07572__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 _01501_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_2
XANTENNA__11218__B top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09313__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__A_N _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ clknet_leaf_48_clk _00510_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07324__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07271__X _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ clknet_leaf_23_clk _00441_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11828_ _05630_ _05655_ _05632_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11759_ _05578_ _05622_ _05623_ _05576_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_43_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload103 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_181_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10284__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ clknet_leaf_4_clk _00993_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06850__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08830__X _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09077__C net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06602__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ _02117_ net591 net1227 net868 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13636__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ top.DUT.register\[20\]\[16\] net748 _03041_ _03047_ vssd1 vssd1 vccd1 vccd1
+ _03048_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_126_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07852_ top.DUT.register\[4\]\[18\] net566 net543 top.DUT.register\[22\]\[18\] _02978_
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a221o_1
XANTENNA__09093__B _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__B _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__inv_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
X_07783_ top.DUT.register\[12\]\[19\] net582 net737 top.DUT.register\[24\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_48_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12206__A2_N _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__A2 _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__A1 _01588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _01797_ _04557_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_211_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06734_ _01840_ _01859_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_203_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07315__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__B net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09453_ _01991_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10459__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06665_ top.DUT.register\[25\]\[27\] net771 net689 top.DUT.register\[3\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout252_A _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ _02516_ _02542_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__nand2_1
X_09384_ _04426_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_135_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06596_ top.DUT.register\[29\]\[29\] net665 net637 top.DUT.register\[16\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08335_ _02683_ net483 net479 _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08266_ net478 _03375_ _03390_ _03256_ _03388_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a221o_2
XANTENNA__07094__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07217_ top.DUT.register\[29\]\[15\] net663 net607 top.DUT.register\[12\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06841__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08197_ _02608_ net294 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nand2_1
XANTENNA__09983__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ net508 _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout886_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _02188_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__nor2_2
XFILLER_0_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10922__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Left_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1007 net1008 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_2
X_10090_ net168 net1773 net418 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1029 net1051 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09571__X _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12800_ clknet_leaf_47_clk _00364_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13780_ clknet_leaf_65_clk _01323_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ top.a1.data\[2\] top.a1.dataInTemp\[6\] net797 vssd1 vssd1 vccd1 vccd1 _05010_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07306__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ clknet_leaf_56_clk _00295_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_153_Left_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12662_ clknet_leaf_121_clk _00226_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _05461_ _05468_ _05449_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_172_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ clknet_leaf_110_clk _00157_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11544_ _05379_ _05407_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06832__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11475_ _05308_ _05323_ net267 _05316_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a31o_1
Xwire498 _02630_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_2
X_13214_ clknet_leaf_13_clk _00778_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ net221 net2011 net325 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_162_Left_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12645__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ clknet_leaf_36_clk _00709_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10832__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357_ net1662 net192 net395 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07793__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13076_ clknet_leaf_60_clk _00640_ net1099 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10288_ net2046 net203 net403 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__mux2_1
X_12027_ _05868_ _05871_ net127 _05872_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_183_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07545__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_171_Left_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12929_ clknet_leaf_27_clk _00493_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10279__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06450_ _01576_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__inv_2
XFILLER_0_201_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06381_ top.a1.instruction\[17\] top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ _01508_ sky130_fd_sc_hd__and2_2
XANTENNA__11899__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08120_ _02143_ net290 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08051_ _03174_ _03175_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_180_Left_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07002_ top.DUT.register\[20\]\[11\] net750 net729 top.DUT.register\[10\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
XANTENNA__09222__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ net1175 net865 _02709_ net593 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_168_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07904_ _03029_ _03030_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_4_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ net280 _03980_ _03981_ net300 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_90_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07904__X _03031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ top.DUT.register\[26\]\[18\] net762 net715 top.DUT.register\[30\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a22o_1
XANTENNA__07000__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ _02516_ _02543_ _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a21o_1
X_09505_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__inv_2
X_06717_ top.DUT.register\[24\]\[26\] net551 net597 top.DUT.register\[27\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10189__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07697_ top.DUT.register\[29\]\[0\] net700 net692 top.DUT.register\[21\]\[0\] _02822_
+ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout634_A _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__B net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ _04444_ _04449_ _04461_ _04462_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__o31a_1
XANTENNA__09978__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06648_ _01755_ _01774_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_109_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09367_ net906 top.pc\[18\] _04403_ _04412_ net896 vssd1 vssd1 vccd1 vccd1 _00099_
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ top.DUT.register\[6\]\[29\] net765 net687 top.DUT.register\[1\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08318_ net302 _03233_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__nand2_1
XANTENNA__09279__A _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08264__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09298_ _04344_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08249_ net283 _03373_ _03368_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06814__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11260_ top.a1.row2\[2\] _05111_ _05100_ _01444_ vssd1 vssd1 vccd1 vccd1 _05138_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ net225 net1825 net406 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__mux2_1
XANTENNA__10652__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ top.a1.row1\[3\] net530 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__and2_1
X_10142_ net232 net1912 net414 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10073_ net235 net2274 net417 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_68_clk _01373_ net1105 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13763_ clknet_leaf_85_clk _01306_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10099__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ top.a1.dataIn\[1\] net848 _04995_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_
+ sky130_fd_sc_hd__a22o_1
X_12714_ clknet_leaf_34_clk _00278_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13694_ clknet_leaf_73_clk _01242_ net1091 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ clknet_leaf_119_clk _00209_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10827__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12576_ clknet_leaf_45_clk _00140_ net1082 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11527_ _05362_ _05383_ _05384_ _05357_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06805__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ _05288_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08821__A _01865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10409_ net160 net2231 net327 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__mux2_1
XANTENNA__10562__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11389_ _01390_ _05256_ _05235_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__a21o_1
X_13128_ clknet_leaf_35_clk _00692_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13059_ clknet_leaf_50_clk _00623_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 top.DUT.register\[24\]\[4\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07518__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09652__A _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ top.DUT.register\[16\]\[2\] net635 net595 top.DUT.register\[27\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09371__B _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_200_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ top.DUT.register\[22\]\[4\] net753 net717 top.DUT.register\[2\]\[4\] _02677_
+ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06502_ top.a1.instruction\[23\] _01627_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_196_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07482_ top.a1.instruction\[25\] _01621_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _04258_ _04260_ _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06433_ _01547_ _01559_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__nor2_8
XANTENNA__10737__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ top.pc\[2\] top.pc\[3\] top.pc\[4\] top.pc\[5\] vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06364_ top.d_ready top.ru.state\[0\] net794 net34 vssd1 vssd1 vccd1 vccd1 _00005_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08103_ _02682_ net295 vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06295_ _01438_ _01439_ _01442_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09083_ _04062_ _04096_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nor3_2
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout215_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ _01569_ _03155_ _03160_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__and3_1
Xhold810 top.DUT.register\[27\]\[9\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 top.DUT.register\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold832 top.DUT.register\[6\]\[22\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 top.DUT.register\[23\]\[0\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11002__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10472__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 top.DUT.register\[15\]\[31\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 top.DUT.register\[29\]\[18\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold876 top.DUT.register\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold887 top.DUT.register\[13\]\[10\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 top.DUT.register\[15\]\[4\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07221__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ net1532 net177 net429 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout584_A _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ net1358 net838 net817 _04031_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__a22o_1
X_08867_ _03889_ _03965_ net305 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__B _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ top.DUT.register\[8\]\[19\] net569 net554 top.DUT.register\[7\]\[19\] _02934_
+ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a221o_1
XANTENNA__08178__A _02143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08798_ _01950_ _03885_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__and2b_1
XANTENNA__06732__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07749_ net494 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10760_ net190 net1731 net375 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__mux2_1
XANTENNA__07288__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09682__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09419_ _02056_ _04460_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or2_1
XANTENNA__10647__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ net230 net1679 net378 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12430_ clknet_leaf_97_clk top.ru.next_FetchedData\[14\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08788__A2 _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12361_ top.pad.button_control.r_counter\[13\] _06144_ vssd1 vssd1 vccd1 vccd1 _06146_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07996__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ top.a1.dataIn\[27\] top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12292_ top.lcd.cnt_500hz\[4\] _01438_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09737__A1 _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ top.a1.row1\[0\] _05094_ _05119_ top.a1.row1\[16\] vssd1 vssd1 vccd1 vccd1
+ _05123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06161__A top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net1463 net532 net525 _05074_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__a22o_1
X_10125_ net1574 net160 net459 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10056_ net170 net2146 net422 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11507__A top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ clknet_leaf_70_clk _01356_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13746_ clknet_leaf_88_clk _01289_ net1006 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07279__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ _04979_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08476__B2 _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13677_ clknet_leaf_94_clk _00005_ net993 vssd1 vssd1 vccd1 vccd1 top.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10557__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10889_ net1703 net203 net347 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12628_ clknet_leaf_47_clk _00192_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__B2 _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ clknet_leaf_20_clk _00123_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09069__D _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09647__A top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07451__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold106 net123 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold117 _01181_ vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold128 top.a1.row1\[121\] vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top.ramaddr\[24\] vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10292__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07739__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07203__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout608 _01667_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout619 _01663_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_186_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06411__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ top.pc\[17\] _04394_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_1
X_06982_ top.DUT.register\[20\]\[20\] net579 net661 top.DUT.register\[2\]\[20\] _02108_
+ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a221o_1
X_08721_ net318 _03447_ _03745_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_198_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09361__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ _03082_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07911__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _02718_ _02719_ _02727_ _02729_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__or4_4
XFILLER_0_95_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08583_ _02402_ net488 net469 _02403_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout165_A _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07534_ net808 _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07465_ top.DUT.register\[26\]\[5\] net759 net708 top.DUT.register\[9\]\[5\] _02591_
+ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10467__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09204_ _04257_ _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nand2_1
XANTENNA__08219__A1 _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06416_ _01496_ net791 _01503_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__and3_4
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08219__B2 _03343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ top.DUT.register\[13\]\[7\] net648 net640 top.DUT.register\[11\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09135_ _01618_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__nand2_1
X_06347_ net903 net901 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__or2_1
XANTENNA__08498__A1_N _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09066_ _02276_ _02318_ _02359_ _02402_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__and4_1
XANTENNA__07442__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06278_ net1635 net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[22\] sky130_fd_sc_hd__and2_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout799_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ top.DUT.register\[7\]\[31\] net554 net625 top.DUT.register\[25\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a22o_1
Xhold640 top.DUT.register\[25\]\[3\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 top.DUT.register\[8\]\[11\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 top.pad.button_control.r_counter\[6\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold673 top.DUT.register\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 top.DUT.register\[21\]\[3\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 top.pad.button_control.r_counter\[5\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ top.DUT.register\[3\]\[6\] net243 net431 vssd1 vssd1 vccd1 vccd1 _00192_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10930__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08919_ net1245 net838 net817 _04015_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09899_ _04891_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11327__A top.a1.dataIn\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11861_ _01398_ net130 _05684_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a21o_1
X_13600_ clknet_leaf_95_clk _01159_ net990 vssd1 vssd1 vccd1 vccd1 top.ramload\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10812_ net1599 net237 net353 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ _05660_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__nor2_1
XANTENNA__08636__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13531_ clknet_leaf_53_clk _01095_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10743_ net252 net1717 net375 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13462_ clknet_leaf_119_clk _01026_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10674_ net1886 net142 net452 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12413_ clknet_leaf_83_clk _00049_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_209_Right_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13393_ clknet_leaf_12_clk _00957_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12344_ _06134_ _06135_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__nor2_1
XANTENNA__09467__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07433__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08371__A _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ _06092_ _06093_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11226_ net891 _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_56_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10840__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ net1293 net533 _05065_ _05066_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ net1616 net226 net459 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11088_ net917 net1301 net852 _05030_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a31o_1
X_10039_ net235 net2245 net421 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
XANTENNA__08697__A1 _03426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08697__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10287__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13729_ clknet_leaf_72_clk _01272_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07250_ top.DUT.register\[24\]\[14\] net737 net672 top.DUT.register\[16\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07672__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06201_ _00009_ top.a1.nextHex\[7\] vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[2\] sky130_fd_sc_hd__or2_1
XANTENNA__06880__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ top.DUT.register\[15\]\[13\] _01655_ net783 top.DUT.register\[31\]\[13\]
+ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08552__Y _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07424__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06632__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout405 _04935_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_6
Xfanout416 _04931_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_4
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_8
X_09822_ _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__nand2_1
XANTENNA__10750__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _04681_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_4
X_09753_ _04751_ _04755_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__and3_1
X_06965_ top.DUT.register\[31\]\[20\] net745 net717 top.DUT.register\[2\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a22o_1
X_08704_ net471 _03798_ _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o21ai_1
X_09684_ _03462_ net340 net336 _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__o211a_2
XANTENNA__08688__A1 _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06896_ top.DUT.register\[24\]\[22\] net550 net601 top.DUT.register\[10\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _03215_ _03240_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__nand2_1
XANTENNA__06699__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ _03620_ _03679_ net280 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__mux2_1
XANTENNA__06528__X _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ top.DUT.register\[3\]\[4\] net787 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10197__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08497_ _03612_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_A _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07448_ top.DUT.register\[20\]\[6\] net579 net598 top.DUT.register\[27\]\[6\] _02574_
+ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07663__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06871__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10925__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07379_ top.DUT.register\[28\]\[7\] net585 net686 top.DUT.register\[1\]\[7\] _02505_
+ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _01406_ _04044_ _04179_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08191__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net238 net1831 net327 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__mux2_1
XANTENNA__07415__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09049_ _03560_ _03579_ _03608_ _03630_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__and4_1
Xclkbuf_4_4__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ _05903_ _05906_ _05922_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a21oi_1
Xhold470 top.DUT.register\[20\]\[22\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold481 top.DUT.register\[25\]\[20\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ net1 wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__nand2_1
Xhold492 top.DUT.register\[26\]\[12\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10660__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net955 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_4
Xfanout961 net964 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_2
Xfanout972 net978 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_2
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ clknet_leaf_43_clk _00526_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1170 top.DUT.register\[20\]\[25\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _05777_ _05779_ _05781_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__and3_1
Xhold1181 top.DUT.register\[7\]\[12\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12893_ clknet_leaf_107_clk _00457_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_206_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11844_ _05705_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11775_ _05643_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08085__B _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13514_ clknet_leaf_38_clk _01078_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10726_ net204 net2042 net384 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08851__B2 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13445_ clknet_leaf_118_clk _01009_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06862__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657_ net2170 net196 net451 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
XANTENNA__10835__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09909__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload15 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_6
Xclkload26 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_4
X_13376_ clknet_leaf_44_clk _00940_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload37 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_6
XANTENNA__07406__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10588_ net231 net2119 net385 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
Xclkload48 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload48/X sky130_fd_sc_hd__clkbuf_8
Xclkload59 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_6
XANTENNA__06614__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12327_ top.pad.button_control.r_counter\[0\] net795 vssd1 vssd1 vccd1 vccd1 _01353_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_39_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08958__A1_N _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_192_Right_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09159__A2 _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ net1737 _06081_ net1107 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_167_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11209_ net1205 net530 _05091_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__a21o_1
XANTENNA__10570__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ net1674 net846 net814 _06057_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06750_ top.DUT.register\[4\]\[25\] net769 net741 top.DUT.register\[8\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a22o_1
XANTENNA__09867__B1 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire515_A _01948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06681_ top.DUT.register\[8\]\[27\] net568 net603 top.DUT.register\[18\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08420_ net482 net275 _03537_ _03525_ net469 vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_69_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13495__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07893__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08351_ _03310_ _03326_ net308 vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07302_ top.DUT.register\[1\]\[9\] net656 net555 top.DUT.register\[7\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a22o_1
X_08282_ _03405_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07645__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__06853__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07233_ _02339_ _02358_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__nor2_1
XANTENNA__10745__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07164_ _02282_ _02283_ _02289_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__or4_4
XFILLER_0_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06605__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07095_ top.DUT.register\[3\]\[10\] net785 _02221_ vssd1 vssd1 vccd1 vccd1 _02222_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_113_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1037_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout202 _04748_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
Xfanout224 _04729_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_1
XANTENNA__09554__B _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07030__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ net834 _04436_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nor2_1
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
Xfanout268 _03187_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
Xfanout279 _02856_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
X_07997_ top.DUT.register\[19\]\[31\] net734 net679 top.DUT.register\[13\]\[31\] _03123_
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06948_ _02065_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nor2_4
X_09736_ net835 _04327_ _04720_ top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 _04746_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08738__X _03844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09667_ top.a1.dataIn\[0\] _01492_ _04689_ top.pc\[0\] net343 vssd1 vssd1 vccd1 vccd1
+ _04690_ sky130_fd_sc_hd__a221o_1
X_06879_ _01999_ _02003_ _02004_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout929_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ net481 _03727_ _03728_ net520 _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__o221a_1
XANTENNA__07802__B net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12209__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ top.a1.state\[2\] net893 top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04630_
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_194_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08549_ _02278_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07097__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11560_ _05385_ _05418_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__xor2_2
XFILLER_0_175_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07636__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__B2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10511_ net147 net1754 net366 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__mux2_1
XANTENNA__06844__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11491_ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__inv_2
XANTENNA__09729__B _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10655__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08633__B net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13230_ clknet_leaf_110_clk _00794_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09389__A2 top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10442_ net160 net1631 net323 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13161_ clknet_leaf_4_clk _00725_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ _01594_ net437 _04687_ net433 vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12112_ _05965_ _05977_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nor2_1
X_13092_ clknet_leaf_40_clk _00656_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10390__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _05906_ _05912_ _05903_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10156__A0 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06440__Y _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07021__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout780 _01682_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_6
Xfanout791 _01501_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__buf_2
XANTENNA__12546__SET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_12_clk _00509_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08096__A _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ clknet_leaf_11_clk _00440_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11827_ _05652_ _05677_ _05691_ _05649_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_190_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07088__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11758_ _05607_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08824__A _01865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10709_ net261 net1931 net381 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XANTENNA__06835__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10565__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11689_ _05552_ _05556_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a31o_2
XFILLER_0_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload104 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_155_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13428_ clknet_leaf_61_clk _00992_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13359_ clknet_leaf_20_clk _00923_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10395__A0 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07260__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ top.DUT.register\[14\]\[16\] net721 net701 top.DUT.register\[29\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a22o_1
XANTENNA__07012__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ top.DUT.register\[23\]\[18\] net563 net553 top.DUT.register\[7\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a22o_1
XANTENNA__07563__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ _01919_ _01928_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__nor2_8
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07782_ _02902_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nand2_1
XANTENNA__09390__A top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A1_N top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ _01797_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06733_ _01840_ _01859_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_211_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ _04303_ _04423_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__and2_1
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06664_ top.DUT.register\[11\]\[27\] net755 net685 top.DUT.register\[1\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08403_ _02516_ _02542_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__or2_2
X_09383_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06595_ top.DUT.register\[8\]\[29\] net569 net625 top.DUT.register\[25\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout245_A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ net321 _03446_ _03442_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07618__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08265_ net313 _03389_ _03364_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a21o_1
XANTENNA__10475__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06525__Y _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07216_ top.DUT.register\[13\]\[15\] net647 net595 top.DUT.register\[27\]\[15\] _02342_
+ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ _03320_ _03321_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07147_ net809 net505 net463 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07251__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06541__X _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ _02192_ _02204_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout781_A _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09284__B _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1019 net1020 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07003__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09719_ top.pc\[11\] net803 _04718_ _04730_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ net1374 _05009_ net535 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__mux2_1
X_12730_ clknet_leaf_19_clk _00294_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07857__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ clknet_leaf_8_clk _00225_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ _05461_ _05469_ _05474_ _05479_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__or4bb_2
XTAP_TAPCELL_ROW_172_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12592_ clknet_leaf_122_clk _00156_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_172_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11543_ top.a1.dataIn\[13\] _05409_ _05410_ _05411_ vssd1 vssd1 vccd1 vccd1 _05413_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06817__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10385__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ _05342_ _05343_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__nor2_1
XANTENNA__07490__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06164__A top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ clknet_leaf_104_clk _00777_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ net225 net1744 net323 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__mux2_1
Xwire499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_2
XFILLER_0_150_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ clknet_leaf_110_clk _00708_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10356_ net1471 net205 net395 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06596__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13075_ clknet_leaf_1_clk _00639_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ net1985 net213 net404 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12026_ _05885_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__or2_1
XANTENNA__11229__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08742__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08538__B net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12928_ clknet_leaf_44_clk _00492_ net1082 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07848__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_52_clk _00423_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06380_ net791 _01505_ _01506_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06808__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10295__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ _03174_ _03175_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__nor2_4
X_07001_ top.DUT.register\[24\]\[11\] net738 net688 top.DUT.register\[1\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06587__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net1354 net865 _02757_ net593 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_168_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ _03014_ _03017_ _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_4_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08883_ net280 _03946_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_205_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout195_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _02954_ _02955_ _02959_ _02960_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__or4_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07765_ _02516_ _02543_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout362_A _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06716_ top.DUT.register\[26\]\[26\] net622 net542 top.DUT.register\[22\]\[26\] _01842_
+ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a221o_1
X_09504_ net528 _04541_ _04423_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07839__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ top.DUT.register\[27\]\[0\] net775 net726 top.DUT.register\[17\]\[0\] _02821_
+ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ net513 _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06647_ net808 net518 net463 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout627_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09366_ net135 _04406_ _04410_ _04411_ net906 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__o221ai_1
XANTENNA__06536__X _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06578_ top.DUT.register\[8\]\[29\] net741 net672 top.DUT.register\[16\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08317_ net303 _03252_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09297_ _04345_ _04346_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__nand2_1
XANTENNA__09279__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08248_ net298 net288 _03127_ _03372_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ net506 net292 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nand2_1
XANTENNA__10933__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08016__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ net231 net1899 net406 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07224__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net1200 net530 _05082_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ net236 top.DUT.register\[8\]\[8\] net413 vssd1 vssd1 vccd1 vccd1 _00354_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ net242 net1580 net417 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
XANTENNA__09921__C1 _04912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13831_ clknet_leaf_68_clk _01372_ net1105 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06750__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13762_ clknet_leaf_85_clk _01305_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10974_ top.a1.halfData\[1\] _04991_ _04996_ net844 vssd1 vssd1 vccd1 vccd1 _04997_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12713_ clknet_leaf_11_clk _00277_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13693_ clknet_leaf_75_clk _01241_ net1090 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ clknet_leaf_33_clk _00208_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ clknet_leaf_115_clk _00139_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11526_ _05368_ _05395_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__and2b_1
XANTENNA__07463__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11457_ _05273_ net331 _05289_ _05290_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08007__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878__1129 vssd1 vssd1 vccd1 vccd1 _13878__1129/HI net1129 sky130_fd_sc_hd__conb_1
XFILLER_0_40_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10408_ net165 net1867 net329 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__mux2_1
XANTENNA__07215__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11388_ _05235_ _05256_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nand2_1
XANTENNA__07766__A1 _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06569__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ net1791 net259 net393 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__mux2_1
X_13127_ clknet_leaf_7_clk _00691_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10770__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ clknet_leaf_43_clk _00622_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12009_ _05849_ net127 vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__and2_1
XANTENNA__09912__C1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06741__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07550_ top.DUT.register\[10\]\[4\] net729 net699 top.DUT.register\[23\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_200_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06501_ top.a1.instruction\[23\] _01627_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07481_ _02599_ _02607_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__nor2_8
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_196_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ top.pc\[9\] _02471_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__xor2_1
X_06432_ _01552_ _01556_ _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__or3_2
XFILLER_0_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ net895 top.pc\[3\] top.pc\[4\] top.pc\[5\] vssd1 vssd1 vccd1 vccd1 _04210_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06363_ _01489_ _01490_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08102_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07454__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ _04115_ _04143_ _04116_ _04105_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_79_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06294_ _01440_ _01441_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08033_ _01570_ _03159_ _02187_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold800 top.DUT.register\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10753__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold811 top.DUT.register\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06803__Y _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__A1 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 top.DUT.register\[2\]\[24\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 top.DUT.register\[24\]\[7\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold844 top.DUT.register\[10\]\[4\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold855 top.DUT.register\[22\]\[0\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 top.DUT.register\[11\]\[11\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__B1 _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 top.DUT.register\[22\]\[2\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 top.DUT.register\[20\]\[20\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 top.DUT.register\[6\]\[6\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net2254 net183 net431 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
X_08935_ net536 _04029_ _04030_ top.pc\[31\] net887 vssd1 vssd1 vccd1 vccd1 _04031_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__06980__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _03928_ _03961_ net277 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__mux2_1
X_07817_ _02936_ _02938_ _02940_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__or4_1
X_08797_ net1299 net839 net817 _03899_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A _01518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06732__A2 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ _02864_ _02867_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nor3_4
XFILLER_0_168_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ top.DUT.register\[21\]\[0\] net572 net627 top.DUT.register\[9\]\[0\] _02805_
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout911_A top.i_ready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10928__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__A1 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09418_ _02056_ _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12573__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ net179 net1813 net377 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
XANTENNA__08194__A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_3__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09434__A1 top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12360_ _06144_ _06145_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__nor2_1
XANTENNA__07445__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11241__B2 top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_X net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06799__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ top.a1.dataIn\[0\] _04629_ net849 _05181_ vssd1 vssd1 vccd1 vccd1 _01274_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12291_ top.lcd.cnt_500hz\[4\] _01438_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or2_1
XANTENNA__10663__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06713__Y _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ top.a1.row1\[120\] _05106_ _05117_ top.a1.row2\[8\] _05121_ vssd1 vssd1 vccd1
+ vccd1 _05122_ sky130_fd_sc_hd__a221o_1
XANTENNA__09737__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11173_ top.a1.dataInTemp\[8\] top.a1.data\[8\] net799 vssd1 vssd1 vccd1 vccd1 _05074_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10752__A0 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ net1808 net166 net460 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ net172 net2260 net423 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07273__A _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08088__B _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06723__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13814_ clknet_leaf_70_clk _01355_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_11_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13745_ clknet_leaf_86_clk _01288_ net1007 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10957_ _01380_ _01418_ _01410_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09673__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10838__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13676_ clknet_leaf_94_clk _00010_ net993 vssd1 vssd1 vccd1 vccd1 top.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10888_ net2293 net213 net348 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ clknet_leaf_1_clk _00191_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__A2 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12558_ clknet_leaf_117_clk _00122_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08832__A _01865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10573__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11509_ top.a1.dataIn\[14\] _05376_ _05377_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__or3_1
XANTENNA__09647__B _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 top.ramstore\[7\] vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ clknet_leaf_114_clk _00056_ net939 vssd1 vssd1 vccd1 vccd1 top.ramstore\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold118 top.DUT.register\[18\]\[15\] vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 top.a1.row1\[113\] vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 _01667_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ top.DUT.register\[17\]\[20\] net646 net559 top.DUT.register\[6\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_165_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_23_clk_X clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _03237_ _03649_ _03825_ net269 _03826_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a221o_1
XANTENNA__09382__B _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08651_ _03035_ _03081_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_198_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ top.DUT.register\[15\]\[3\] net704 net674 top.DUT.register\[18\]\[3\] _02728_
+ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net320 _03694_ _03693_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ _02646_ _02657_ _02658_ _02659_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__or4_4
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10748__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_A _04890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07675__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ top.DUT.register\[27\]\[5\] net775 net772 top.DUT.register\[25\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06415_ top.DUT.register\[29\]\[30\] net701 net690 top.DUT.register\[3\]\[30\] _01534_
+ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__a221o_1
X_09203_ top.pc\[8\] _02521_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08219__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07395_ top.DUT.register\[3\]\[7\] net786 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout325_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _04159_ _04163_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__a21o_1
XANTENNA__07427__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06346_ top.a1.instruction\[6\] _01477_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_146_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09065_ _02163_ _02949_ _02992_ _03033_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__and4_1
XANTENNA__10483__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06277_ top.ramload\[21\] net878 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08016_ top.DUT.register\[11\]\[31\] net641 net628 top.DUT.register\[9\]\[31\] _03131_
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a221o_1
XANTENNA__09719__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 top.DUT.register\[6\]\[19\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 top.DUT.register\[12\]\[7\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 top.DUT.register\[17\]\[30\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold663 top.DUT.register\[4\]\[4\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 top.DUT.register\[9\]\[31\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 top.DUT.register\[17\]\[24\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 top.DUT.register\[31\]\[15\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_A _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ net1439 net246 net429 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__Y _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net887 top.pc\[30\] net536 _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a22o_1
X_09898_ top.pc\[29\] _04587_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__or2_1
XANTENNA__09860__X _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ net318 _03625_ _03804_ _03237_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a221o_2
XANTENNA__06705__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ top.a1.dataIn\[5\] _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13877__1128 vssd1 vssd1 vccd1 vccd1 _13877__1128/HI net1128 sky130_fd_sc_hd__conb_1
XFILLER_0_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ net1579 net242 net354 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__mux2_1
X_11791_ _05633_ _05659_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__and2_1
XANTENNA__10658__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07666__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ clknet_leaf_15_clk _01094_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10742_ net255 net2154 net373 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07130__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09407__A1 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13461_ clknet_leaf_8_clk _01025_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10673_ net2152 net147 net453 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07418__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ clknet_leaf_84_clk _00048_ net1014 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13392_ clknet_leaf_0_clk _00956_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12343_ net1822 _06132_ net796 vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10393__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06206__A_N top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12274_ net2031 _06091_ net1107 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08918__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ net881 _05096_ _05101_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__and3_2
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07197__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ top.a1.data\[0\] net798 _04992_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__o21a_1
XANTENNA__06944__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ net1418 net234 net461 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07274__Y _02401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ net65 net861 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__and2_1
X_10038_ net240 net2300 net421 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08697__A2 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10568__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _05858_ _05799_ _05850_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13728_ clknet_leaf_72_clk _01271_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06347__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08854__C1 _03953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13659_ clknet_leaf_75_clk _01218_ net1017 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06200_ _01424_ net1472 _01419_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[1\] sky130_fd_sc_hd__mux2_1
XANTENNA__07409__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ top.DUT.register\[19\]\[13\] net633 net787 top.DUT.register\[3\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08909__B1 _03878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout406 _04935_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_4
Xfanout417 _04927_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_6
X_09821_ top.pc\[22\] _04476_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__or2_1
XANTENNA__09393__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07906__A _03012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout428 _04923_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_8
Xfanout439 _04681_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_6
XANTENNA__06935__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__A top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ top.pc\[15\] _04362_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__xnor2_1
X_06964_ top.DUT.register\[24\]\[20\] net737 _01535_ top.DUT.register\[3\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22o_1
XANTENNA__08137__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09334__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ net520 _03799_ _03807_ net482 _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__o221a_1
XANTENNA__11147__B _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06895_ top.DUT.register\[9\]\[22\] net629 net610 top.DUT.register\[12\]\[22\] _02021_
+ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a221o_1
X_09683_ net344 _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ net313 _03127_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__nand2_2
XANTENNA__07896__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07360__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08565_ _03301_ _03305_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10478__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07516_ top.DUT.register\[9\]\[4\] net628 net601 top.DUT.register\[10\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ _02235_ _03611_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07112__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07447_ top.DUT.register\[25\]\[6\] net626 net601 top.DUT.register\[10\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11313__D top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A _01533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06544__X _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ top.DUT.register\[26\]\[7\] net759 net726 top.DUT.register\[17\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06329_ _01332_ _01460_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__nand2_1
X_09117_ net895 _04166_ _04177_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ net319 _03628_ _04107_ _04108_ _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__06379__A_N top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold460 top.DUT.register\[5\]\[0\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08972__A2_N net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold471 top.DUT.register\[16\]\[27\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 top.DUT.register\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net918 _01401_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__nor2_1
XANTENNA__07179__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 top.DUT.register\[7\]\[25\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10513__Y _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06926__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net980 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_2
Xfanout951 net954 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
Xfanout962 net964 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12973__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout973 net978 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
Xfanout984 net986 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_129_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ clknet_leaf_28_clk _00525_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1160 top.DUT.register\[18\]\[22\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1171 top.DUT.register\[20\]\[30\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 top.ramload\[5\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _05779_ _05781_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__and2_1
XANTENNA__07887__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 top.ramload\[5\] vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12892_ clknet_leaf_55_clk _00456_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_206_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07351__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10388__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11843_ _05705_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_197_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09628__A1 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07639__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ _01396_ _05638_ _05619_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06167__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ clknet_leaf_3_clk _01077_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ net212 net2296 net384 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
XANTENNA__08653__Y _03763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13444_ clknet_leaf_39_clk _01008_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10656_ net1377 net199 net451 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_12
XFILLER_0_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13375_ clknet_leaf_113_clk _00939_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10587_ net235 net2349 net385 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
Xclkload27 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_8
XFILLER_0_180_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload38 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinv_16
XANTENNA__09800__A1 top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload49 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload49/X sky130_fd_sc_hd__clkbuf_4
X_12326_ _04036_ _04037_ _06122_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__o211a_1
XANTENNA__07811__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ top.lcd.cnt_20ms\[8\] _06081_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__and2_1
XANTENNA__10851__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08367__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08367__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11208_ net850 _05077_ net531 vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__and3_1
X_12188_ _06046_ _06054_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06917__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11139_ net61 net858 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07590__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12605__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07878__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ top.DUT.register\[2\]\[27\] net659 net556 top.DUT.register\[6\]\[27\] _01806_
+ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a221o_1
XFILLER_0_203_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire508_A _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06550__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ net308 _03303_ _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08281_ _03403_ _03404_ net308 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11270__X _05147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07232_ _02339_ _02358_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__and2_2
XFILLER_0_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07163_ top.DUT.register\[19\]\[13\] net733 net730 top.DUT.register\[10\]\[13\] _02286_
+ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06605__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__X _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ top.DUT.register\[31\]\[10\] net781 net779 top.DUT.register\[15\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13876__1127 vssd1 vssd1 vccd1 vccd1 _13876__1127/HI net1127 sky130_fd_sc_hd__conb_1
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10761__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout203 net206 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
Xfanout214 _04795_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout392_A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _04729_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
Xfanout236 net238 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
Xfanout247 net249 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
X_09804_ _04803_ _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__xnor2_1
Xfanout258 _04699_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 _03187_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
X_07996_ top.DUT.register\[6\]\[31\] net765 net718 top.DUT.register\[2\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a22o_1
XANTENNA__07581__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ net823 _01613_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__nor2_1
X_06947_ _02067_ _02069_ _02071_ _02073_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__or4_1
XANTENNA__09858__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07869__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ net534 _04151_ _04682_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__o21a_1
X_06878_ top.DUT.register\[11\]\[22\] net758 net737 top.DUT.register\[24\]\[22\] _01997_
+ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a221o_1
XANTENNA__08467__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__X _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _02360_ net486 net470 _02361_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a22oi_2
XANTENNA_fanout824_A _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ _01384_ top.a1.halfData\[3\] _01385_ _01412_ vssd1 vssd1 vccd1 vccd1 _04629_
+ sky130_fd_sc_hd__or4b_4
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09997__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08548_ _03612_ _03662_ _02163_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08479_ _02235_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__xor2_1
XANTENNA__08833__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ net154 net2171 net367 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__mux2_1
X_11490_ _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10441_ net166 net1298 net325 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06434__B net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__B1 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ clknet_leaf_35_clk _00724_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10372_ net466 _04932_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__nand2_4
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ _05967_ _05975_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10671__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ clknet_leaf_33_clk _00655_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12042_ _05911_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__inv_2
Xhold290 top.DUT.register\[14\]\[23\] vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07572__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout770 _01507_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_4
Xfanout781 _01659_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
Xfanout792 _01500_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_4
X_12944_ clknet_leaf_122_clk _00508_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08521__B2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12875_ clknet_leaf_30_clk _00439_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _05652_ _05677_ _05691_ _05649_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a22oi_2
XANTENNA__08809__C1 _03910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09700__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11757_ _05547_ _05567_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__nand2_1
XANTENNA__10846__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__A2_N net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10708_ net263 net2130 net384 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XANTENNA__08316__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _05496_ _05554_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload105 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__clkinv_4
X_13427_ clknet_leaf_4_clk _00991_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11250__B _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ net156 net1967 net392 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_117_clk _00922_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_188_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12309_ _06113_ net588 _06112_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__and3b_1
XANTENNA__10581__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07727__Y _02854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13289_ clknet_leaf_4_clk _00853_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire458_A _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07850_ top.DUT.register\[28\]\[18\] net654 net610 top.DUT.register\[12\]\[18\] _02976_
+ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_3_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06801_ _01920_ _01923_ _01925_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__or4_4
XFILLER_0_127_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07781_ _02497_ _02893_ _02907_ _02404_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__o22a_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
XANTENNA__06771__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07462__Y _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ net528 _04556_ _04423_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__o21a_2
X_06732_ net806 _01858_ _01624_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_84_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07191__A _02298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _02015_ _04476_ _04479_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a21oi_1
X_06663_ _01782_ _01783_ _01788_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__or4_2
XFILLER_0_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08402_ net1330 net837 net816 _03522_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09382_ _04425_ _02928_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__and2b_1
X_06594_ top.DUT.register\[17\]\[29\] net645 net609 top.DUT.register\[12\]\[29\] _01720_
+ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _03185_ _03455_ net304 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__mux2_2
XFILLER_0_176_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10756__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout140_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ net283 _03372_ _03368_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a21o_1
XANTENNA__11280__C1 _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07215_ top.DUT.register\[11\]\[15\] net639 net611 top.DUT.register\[14\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08195_ net499 net290 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nand2_1
XANTENNA__09225__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_A _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09846__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _02257_ _02259_ _02271_ _02272_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__nor4_1
XFILLER_0_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07077_ _02198_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__nor2_1
XANTENNA__10491__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07366__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 net1019 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XANTENNA__12527__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_A _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_X net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _01733_ _03104_ _01694_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_126_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11175__X _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__A top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ net835 _04295_ _04720_ top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 _04730_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08197__A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ top.a1.dataIn\[5\] net848 net843 _05008_ vssd1 vssd1 vccd1 vccd1 _05009_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07306__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11102__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _01618_ _04158_ _04672_ _04625_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12660_ clknet_leaf_60_clk _00224_ net1102 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11611_ _05461_ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10666__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12591_ clknet_leaf_50_clk _00155_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_67_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _05410_ _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11271__C1 _05147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06445__A top.a1.instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_208_Left_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11473_ _05325_ _05326_ net267 vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__and3_1
Xwire467 _02830_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_137_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13212_ clknet_leaf_17_clk _00776_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10424_ net232 net1417 net324 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08660__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11574__B1 top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_107_clk _00707_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ net1728 net211 net395 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07793__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13074_ clknet_leaf_52_clk _00638_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10286_ net2201 net216 net401 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_76_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12025_ _05860_ _05861_ net127 _05864_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_183_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07545__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06753__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12927_ clknet_leaf_114_clk _00491_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13875__1126 vssd1 vssd1 vccd1 vccd1 _13875__1126/HI net1126 sky130_fd_sc_hd__conb_1
XFILLER_0_158_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12858_ clknet_leaf_18_clk _00422_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_85_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06907__X _02034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _05641_ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10576__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_107_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12789_ clknet_leaf_5_clk _00353_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07000_ top.DUT.register\[3\]\[11\] net691 net679 top.DUT.register\[13\]\[11\] _02124_
+ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ net1307 net868 _02854_ net593 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_168_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07902_ _03022_ _03023_ _03025_ _03028_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__or4_1
X_08882_ _03282_ _03290_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09930__A0 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__A2 _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07833_ top.DUT.register\[10\]\[18\] net729 net723 top.DUT.register\[14\]\[18\] _02956_
+ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07764_ _02562_ _02586_ _02890_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09503_ top.a1.instruction\[26\] net822 _04540_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__o21a_1
X_06715_ top.DUT.register\[7\]\[26\] net553 net629 top.DUT.register\[9\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
X_07695_ top.DUT.register\[24\]\[0\] net735 net696 top.DUT.register\[23\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout355_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1097_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ top.a1.instruction\[22\] net821 _02208_ _04424_ vssd1 vssd1 vccd1 vccd1 _04476_
+ sky130_fd_sc_hd__o31a_2
X_06646_ _01768_ _01770_ _01772_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_121_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09365_ _04408_ _04409_ _01618_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10486__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_A _03183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ _01697_ _01698_ _01702_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__or4_4
XFILLER_0_176_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08316_ _03218_ _03245_ net303 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09296_ top.pc\[14\] _04329_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nand2_1
XANTENNA__09279__C _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ net302 _03371_ _03370_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09576__A _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08178_ _02143_ net297 vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout891_A top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09295__B _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ top.DUT.register\[14\]\[12\] net614 net608 top.DUT.register\[12\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ net239 net1914 net413 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__mux2_1
XANTENNA__11308__B1 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _04711_ net2059 net420 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__B2 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10531__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13830_ clknet_leaf_68_clk _01371_ net1104 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08488__A0 _03386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13761_ clknet_leaf_74_clk _01304_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10973_ top.a1.dataInTemp\[1\] net800 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ clknet_leaf_31_clk _00276_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ clknet_leaf_73_clk _01240_ net1094 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07160__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12643_ clknet_leaf_41_clk _00207_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10396__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11081__A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ clknet_leaf_13_clk _00138_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ _05366_ _05391_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_152_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08661__Y _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09486__A top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _05279_ _05312_ _05309_ net331 vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ net169 net2276 net328 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__mux2_1
X_11387_ _01390_ _05256_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_185_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07766__A2 _02543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ clknet_leaf_24_clk _00690_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08963__B2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10338_ net1494 net265 net395 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__mux2_1
XANTENNA__06974__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ clknet_leaf_25_clk _00621_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ net1501 net150 net401 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07518__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _05856_ _05874_ _05876_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_187_Right_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06500_ top.a1.instruction\[22\] net801 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ _02600_ _02602_ _02604_ _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__or4_4
XFILLER_0_124_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_196_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06431_ top.DUT.register\[26\]\[30\] net760 net713 top.DUT.register\[30\]\[30\] _01557_
+ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06362_ net902 _01479_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__nand2_1
X_09150_ net908 top.pc\[4\] _04209_ net898 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12144__A_N top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08101_ _02516_ net289 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__nand2_1
X_06293_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\] top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__or4b_1
XFILLER_0_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09081_ _04117_ _04122_ _04123_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_79_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09396__A top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ _01581_ _01595_ _03157_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold801 top.DUT.register\[3\]\[25\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 top.DUT.register\[11\]\[10\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 top.DUT.register\[19\]\[17\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11002__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold834 top.a1.row1\[108\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold845 top.DUT.register\[12\]\[12\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold856 top.DUT.register\[11\]\[25\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 top.DUT.register\[18\]\[5\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 top.DUT.register\[30\]\[13\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08954__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ net2006 net190 net431 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
Xhold889 top.DUT.register\[25\]\[10\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ _04012_ _04028_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ net315 _03657_ _03543_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o21a_1
XANTENNA__06717__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout472_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ top.DUT.register\[30\]\[19\] net617 net609 top.DUT.register\[12\]\[19\] _02942_
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08796_ net886 top.pc\[24\] net536 _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07747_ _02869_ _02871_ _02873_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__or3_1
XANTENNA__09667__C1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11316__D top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07678_ top.DUT.register\[13\]\[0\] net647 net607 top.DUT.register\[12\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a22o_1
XANTENNA__09682__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09417_ net821 _02424_ _04424_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06629_ top.DUT.register\[25\]\[28\] net625 net597 top.DUT.register\[27\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout904_A top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__B1 _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ _03002_ _03011_ _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_101_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09279_ _02291_ _02297_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or3_2
XFILLER_0_118_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07996__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ top.a1.row2\[0\] net847 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__and2_1
X_12290_ _01438_ net588 _06101_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_134_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11241_ top.a1.row2\[0\] _05111_ _05113_ top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1
+ _05121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06442__B _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11172_ net1878 net533 _04636_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__a21o_1
XANTENNA__06956__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ net1653 net170 net461 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ net176 net1668 net421 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__mux2_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06708__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07381__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13813_ clknet_leaf_70_clk net1232 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07920__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13330__RESET_B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13744_ clknet_leaf_86_clk _01287_ net1016 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10956_ _01410_ _04979_ _04983_ _04984_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__a31o_1
XANTENNA__07133__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07684__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13675_ clknet_leaf_92_clk _01233_ net1000 vssd1 vssd1 vccd1 vccd1 top.busy_o sky130_fd_sc_hd__dfrtp_4
X_10887_ top.DUT.register\[30\]\[17\] net216 net345 vssd1 vssd1 vccd1 vccd1 _01067_
+ sky130_fd_sc_hd__mux2_1
X_12626_ clknet_leaf_49_clk _00190_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09768__X _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_159_Left_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09425__A2 top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07436__A1 top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07436__B2 top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10854__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ clknet_leaf_103_clk _00121_ net1001 vssd1 vssd1 vccd1 vccd1 top.pc\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09830__C1 _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08832__B _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07729__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ _05376_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__or2_1
XANTENNA__07987__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ clknet_leaf_75_clk _00055_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold108 _01174_ vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 top.ramaddr\[22\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ _05289_ _05290_ _05272_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12193__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07739__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13109_ clknet_leaf_6_clk _00673_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06411__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06980_ top.DUT.register\[26\]\[20\] net621 net543 top.DUT.register\[22\]\[20\] _02106_
+ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_168_Left_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08650_ _03035_ _03759_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07372__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ top.DUT.register\[4\]\[3\] net767 net708 top.DUT.register\[9\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XANTENNA__07911__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ net283 _03495_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__or2_2
XFILLER_0_135_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11714__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ top.DUT.register\[8\]\[4\] net569 net542 top.DUT.register\[22\]\[4\] _02647_
+ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07463_ top.DUT.register\[29\]\[5\] net700 net692 top.DUT.register\[21\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ _02521_ top.pc\[8\] vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nand2b_1
X_06414_ _01496_ _01497_ net790 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ top.a1.instruction\[28\] net528 _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_134_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _04192_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__nand2_1
X_06345_ _01475_ net905 net904 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10764__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout220_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06276_ net2156 net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[20\] sky130_fd_sc_hd__and2_1
X_09064_ _01952_ _02234_ net487 _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08015_ top.DUT.register\[4\]\[31\] net566 net542 top.DUT.register\[22\]\[31\] _03130_
+ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_116_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold620 top.DUT.register\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 top.DUT.register\[14\]\[2\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 top.DUT.register\[19\]\[5\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12184__B1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold653 top.DUT.register\[24\]\[15\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09854__A top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 top.DUT.register\[15\]\[3\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 top.DUT.register\[22\]\[29\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 top.DUT.register\[19\]\[11\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 top.DUT.register\[12\]\[9\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ net1816 net254 net431 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
XANTENNA__09573__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _04012_ _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__nor2_1
X_09897_ top.pc\[29\] _04587_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_96_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ net300 _03947_ _03945_ net269 vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07661__X _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ net890 top.pc\[23\] net539 _03882_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a22o_1
XANTENNA__12204__A2_N _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ top.DUT.register\[28\]\[6\] net245 net356 vssd1 vssd1 vccd1 vccd1 _00992_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ _05633_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__nor2_1
XANTENNA__07115__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ net261 net2263 net373 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ clknet_leaf_62_clk _01024_ net1102 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10672_ top.DUT.register\[23\]\[29\] net152 net451 vssd1 vssd1 vccd1 vccd1 _00855_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ clknet_leaf_86_clk _00047_ net1014 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13391_ clknet_leaf_22_clk _00955_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10674__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12342_ top.pad.button_control.r_counter\[6\] _06132_ vssd1 vssd1 vccd1 vccd1 _06134_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06453__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ top.lcd.cnt_20ms\[14\] _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11224_ net884 _05095_ _05101_ net882 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__and4b_1
XFILLER_0_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07555__Y _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ top.a1.state\[2\] net533 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10106_ net2217 net235 net459 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11086_ net915 net1376 net853 _05029_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_147_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08099__B _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10037_ net244 net1632 net423 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
XANTENNA__07354__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10849__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11988_ _05800_ _05832_ _05829_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13727_ clknet_leaf_72_clk _01270_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfxtp_1
X_10939_ net912 _04967_ net798 net843 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13658_ clknet_leaf_83_clk _01217_ net1013 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_30_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08843__A _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12609_ clknet_leaf_28_clk _00173_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06880__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10584__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11205__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ clknet_leaf_98_clk _01148_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06363__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06632__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09820_ top.pc\[22\] _04476_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nand2_1
XANTENNA__09582__A1 _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 _04935_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_6
Xfanout418 _04927_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_4
Xfanout429 _04920_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07593__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _04362_ net527 _04758_ _04718_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a211o_1
X_06963_ top.DUT.register\[4\]\[20\] net768 net707 top.DUT.register\[15\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_78_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09334__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ _03431_ _03771_ _03809_ _02949_ _03808_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o221a_1
X_09682_ top.a1.dataIn\[4\] net794 net803 top.pc\[4\] _04700_ vssd1 vssd1 vccd1 vccd1
+ _04701_ sky130_fd_sc_hd__a221o_1
X_06894_ top.DUT.register\[29\]\[22\] net665 net642 top.DUT.register\[11\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
X_08633_ net321 net490 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nor2_1
XANTENNA__06699__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10759__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08564_ net320 _03677_ _03674_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__o21a_1
X_07515_ _02641_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08495_ _02235_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07446_ top.DUT.register\[21\]\[6\] net574 net543 top.DUT.register\[22\]\[6\] _02572_
+ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10494__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ top.DUT.register\[20\]\[7\] net747 net711 top.DUT.register\[9\]\[7\] _02503_
+ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout602_A _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ net910 net897 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__nand2_2
X_06328_ _01332_ _01463_ _01467_ _01450_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
XANTENNA__08073__A1 _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09270__B1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10955__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06623__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ net313 _03654_ _04088_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06259_ net1359 net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[3\] sky130_fd_sc_hd__and2_1
XANTENNA__09022__B1 _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 top.DUT.register\[30\]\[4\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold461 top.DUT.register\[31\]\[18\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 top.DUT.register\[5\]\[6\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold483 top.DUT.register\[18\]\[4\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 top.DUT.register\[4\]\[22\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07584__A0 _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net933 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09871__X _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout941 net946 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_4
X_09949_ net189 top.DUT.register\[2\]\[21\] net435 vssd1 vssd1 vccd1 vccd1 _00175_
+ sky130_fd_sc_hd__mux2_1
Xfanout952 net954 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 net964 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_205_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net978 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
Xfanout985 net986 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ clknet_leaf_44_clk _00524_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1150 top.DUT.register\[10\]\[24\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ _05722_ _05723_ _05780_ _05758_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__a31o_1
Xhold1161 net72 vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 top.DUT.register\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1183 top.DUT.register\[29\]\[4\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10669__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ clknet_leaf_52_clk _00455_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1194 top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
X_11842_ _05671_ _05709_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_142_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06448__A top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11773_ _01396_ _05619_ _05638_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ clknet_leaf_35_clk _01076_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ net215 net2044 net381 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13443_ clknet_leaf_33_clk _01007_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06862__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ net1505 net208 net451 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
XANTENNA__12185__A top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload17 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_8
X_13374_ clknet_leaf_12_clk _00938_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload28 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload28/X sky130_fd_sc_hd__clkbuf_8
X_10586_ net239 net2210 net386 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
XANTENNA__09800__A2 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload39 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_58_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12325_ top.pad.button_control.debounce top.pad.button_control.noisy vssd1 vssd1
+ vccd1 vccd1 _06123_ sky130_fd_sc_hd__nand2_1
XANTENNA__06614__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12256_ _06081_ net1108 _06080_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_71_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ net1197 net530 _05090_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__a21o_1
X_12187_ net1326 net846 net814 _06056_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07575__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11138_ net917 net1247 net852 _05055_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__a31o_1
XANTENNA__12421__Q top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ net85 net863 net826 net1227 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07327__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_clk_X clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07300_ top.a1.instruction\[30\] net529 _02426_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13423__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08280_ _03270_ _03274_ net282 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07231_ net809 net504 net463 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06853__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07162_ top.DUT.register\[12\]\[13\] net583 net722 top.DUT.register\[14\]\[13\] _02287_
+ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07093_ top.DUT.register\[1\]\[10\] net656 net552 top.DUT.register\[7\]\[10\] _02219_
+ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a221o_1
XANTENNA__06605__A2 _01731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13433__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout204 net206 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06369__A1 top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout215 net218 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07566__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _04729_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_1
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_2
X_09803_ _04804_ _04805_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07030__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
Xfanout259 net262 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
X_07995_ top.DUT.register\[22\]\[31\] net753 net683 top.DUT.register\[7\]\[31\] _03121_
+ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout385_A _04945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _04742_ _04743_ net802 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__and3b_1
X_06946_ top.DUT.register\[28\]\[21\] net654 net565 top.DUT.register\[4\]\[21\] _02072_
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a221o_1
XANTENNA__11114__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ net34 _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__and2_1
X_06877_ top.DUT.register\[12\]\[22\] net583 net679 top.DUT.register\[13\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout552_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08616_ _03543_ _03718_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__nand2_1
X_09596_ top.a1.halfData\[3\] top.a1.halfData\[0\] _01412_ top.a1.halfData\[5\] vssd1
+ vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__and4b_1
X_08547_ _02164_ _02233_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07097__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A1 _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06555__X _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ _02903_ _03574_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07429_ top.DUT.register\[26\]\[6\] net762 net699 top.DUT.register\[23\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a22o_1
XANTENNA__06844__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10440_ net170 net1710 net324 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ _01601_ net465 _04921_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__nor3_1
XFILLER_0_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _05971_ _05975_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__or2_1
X_13090_ clknet_leaf_43_clk _00654_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12041_ _05904_ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 top.DUT.register\[13\]\[8\] vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 top.DUT.register\[27\]\[26\] vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07021__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 _01510_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout771 _01504_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_6
Xfanout782 _01659_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout793 _01500_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12943_ clknet_leaf_20_clk _00507_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10399__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ clknet_leaf_38_clk _00438_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _05689_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__nand2_1
XANTENNA__08809__B1 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ _05621_ _05624_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__and3_1
XANTENNA__07088__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ net148 net1253 net381 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06835__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ _05494_ _05542_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13426_ clknet_leaf_51_clk _00990_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10638_ net160 net2101 net389 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__mux2_1
XANTENNA__11250__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload106 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12416__Q top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10862__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_32_clk _00921_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10569_ net183 net1630 net359 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07796__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ top.lcd.cnt_500hz\[9\] top.lcd.cnt_500hz\[10\] _06109_ vssd1 vssd1 vccd1
+ vccd1 _06113_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_188_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13288_ clknet_leaf_35_clk _00852_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07260__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ _01383_ _06071_ net1107 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o21a_1
XANTENNA__07548__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07012__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06800_ top.DUT.register\[15\]\[24\] net706 net683 top.DUT.register\[7\]\[24\] _01926_
+ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a221o_1
XANTENNA__08760__A2 top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ _02279_ _02903_ _02906_ _02277_ _02904_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__o221a_1
XANTENNA__08568__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
X_06731_ _01843_ _01855_ _01856_ _01857_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__or4_4
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ _04488_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__xnor2_1
X_06662_ top.DUT.register\[12\]\[27\] net580 net700 top.DUT.register\[29\]\[27\] _01786_
+ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a221o_1
XANTENNA__10102__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__A_N _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__X _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08401_ net887 top.pc\[6\] net538 _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a22o_1
XANTENNA__12813__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09381_ _02928_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__nand2b_1
X_06593_ top.DUT.register\[21\]\[29\] net575 net653 top.DUT.register\[28\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08971__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ _03384_ _03454_ net277 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06375__X _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08263_ net473 _03377_ _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout133_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07214_ top.DUT.register\[17\]\[15\] net643 net556 top.DUT.register\[6\]\[15\] _02340_
+ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08194_ _02516_ net295 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ top.DUT.register\[24\]\[12\] net550 net547 top.DUT.register\[5\]\[12\] _02260_
+ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07787__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07076_ _01481_ _01571_ _02199_ _02202_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__o211a_1
XANTENNA__07251__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09528__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__B _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07003__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08749__Y _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07653__Y _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ _01733_ _03104_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09717_ net223 top.DUT.register\[1\]\[10\] net438 vssd1 vssd1 vccd1 vccd1 _00132_
+ sky130_fd_sc_hd__mux2_1
X_06929_ _02045_ _02050_ _02055_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__or3_4
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _04156_ _04157_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__or2_1
XANTENNA__10012__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07711__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _04611_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11610_ _05474_ _05479_ _05469_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12590_ clknet_leaf_117_clk _00154_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08267__B2 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11541_ _01393_ net250 _05378_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_122_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06817__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06445__B top.a1.instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11472_ _05325_ _05331_ _05326_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07490__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ clknet_leaf_59_clk _00775_ net1109 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10423_ net237 net2065 net323 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__mux2_1
XANTENNA__09767__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10682__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06732__Y _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07557__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ clknet_leaf_2_clk _00706_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10354_ net1606 net217 net393 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07242__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__A1 top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ clknet_leaf_12_clk _00637_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10285_ net1672 net229 net402 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
X_12024_ _05891_ _05892_ _05884_ _05889_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_131_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08742__A2 top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07563__Y _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _06060_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_205_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06179__Y _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ clknet_leaf_15_clk _00490_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10857__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ clknet_leaf_36_clk _00421_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08137__B1_N net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ _05672_ _05676_ _05646_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_140_Left_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12788_ clknet_leaf_60_clk _00352_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09012__A _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11739_ _05514_ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06808__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10592__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__B2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_27_clk _00973_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08950_ net1214 net867 _02808_ net593 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__a22o_1
X_07901_ top.DUT.register\[5\]\[17\] net544 net611 top.DUT.register\[14\]\[17\] _03027_
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_168_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ _01736_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_4_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08569__Y _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ top.DUT.register\[4\]\[18\] net769 net587 top.DUT.register\[28\]\[18\] _02957_
+ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_90_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12660__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ _02589_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09502_ _01564_ _02734_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__or2_1
X_06714_ top.DUT.register\[19\]\[26\] net633 net787 top.DUT.register\[3\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07694_ top.DUT.register\[31\]\[0\] net743 net708 top.DUT.register\[9\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a22o_1
XANTENNA__11096__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09694__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ _04471_ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06645_ top.DUT.register\[28\]\[28\] net654 net553 top.DUT.register\[7\]\[28\] _01771_
+ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10767__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout348_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _04408_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08237__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06576_ top.DUT.register\[11\]\[29\] net757 net737 top.DUT.register\[24\]\[29\] _01700_
+ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a221o_1
X_08315_ net1301 net839 net815 _03438_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09295_ top.pc\[14\] _04329_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ net288 _03202_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11005__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06680__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ net280 _03301_ _03302_ _03300_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a31o_1
XANTENNA__12709__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12283__A _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07128_ net507 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__inv_2
XANTENNA__07224__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07059_ top.a1.instruction\[20\] net524 _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a21o_1
XANTENNA__10007__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10070_ net246 net1980 net417 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09921__A1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__B2 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13760_ clknet_leaf_74_clk _01303_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10972_ top.a1.halfData\[1\] net798 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__or2_1
X_12711_ clknet_leaf_8_clk _00275_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10677__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13691_ clknet_leaf_75_clk _01239_ net1090 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ clknet_leaf_41_clk _00206_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11081__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__B1 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12573_ clknet_leaf_104_clk _00137_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11524_ _05390_ _05393_ _05389_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07463__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06671__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__Y _02685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ _05301_ _05307_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ net172 net1977 net330 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07215__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11386_ _05248_ _05254_ _05255_ _05223_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13125_ clknet_leaf_116_clk _00689_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06423__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ net1935 net148 net393 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13056_ clknet_leaf_44_clk _00620_ net1082 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ net466 _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__nor2_4
XFILLER_0_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09912__A1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ _05856_ _05874_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09912__B2 top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ _04916_ _04929_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__nor2_2
XANTENNA__07923__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07750__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10587__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12909_ clknet_leaf_23_clk _00473_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13889_ net1139 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_196_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06430_ top.DUT.register\[6\]\[30\] net764 net736 top.DUT.register\[24\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13277__RESET_B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06361_ net902 _01479_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__and2_1
X_08100_ _02562_ net295 vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09080_ _04130_ _04135_ _04141_ _02497_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__o22ai_1
X_06292_ top.lcd.cnt_500hz\[8\] top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\] top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__or4b_1
XANTENNA__07454__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_204_Right_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08031_ net901 _01577_ _01578_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__or3_1
XFILLER_0_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06662__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09396__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold802 top.DUT.register\[10\]\[21\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold813 top.DUT.register\[26\]\[6\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07206__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold824 top.a1.data\[2\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold835 top.DUT.register\[22\]\[25\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 top.DUT.register\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 top.DUT.register\[12\]\[23\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08954__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ top.DUT.register\[3\]\[20\] net191 net432 vssd1 vssd1 vccd1 vccd1 _00206_
+ sky130_fd_sc_hd__mux2_1
Xhold868 top.DUT.register\[5\]\[21\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 top.DUT.register\[6\]\[21\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ _04012_ _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09903__A1 _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__A2 top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _01776_ net485 _03962_ _01777_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07914__B1 _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07952__A_N _03012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ top.DUT.register\[11\]\[19\] net641 net784 top.DUT.register\[31\]\[19\] _02941_
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a221o_1
X_08795_ _03331_ _03886_ _03895_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a211oi_4
X_07746_ top.DUT.register\[29\]\[1\] net702 net676 top.DUT.register\[18\]\[1\] _02872_
+ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a221o_1
XANTENNA__09667__B1 _04689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13507__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _02796_ _02798_ _02800_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__or4_1
XANTENNA__10497__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout632_A _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09416_ _04444_ _04449_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nor2_1
X_06628_ _01749_ _01754_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__nor2_8
XFILLER_0_137_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09347_ _01615_ _02563_ _02610_ net821 _01622_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__o221a_2
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06559_ _01677_ _01679_ _01681_ _01685_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_101_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07445__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ _01615_ _02736_ _02786_ net823 _01622_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__o221a_4
XTAP_TAPCELL_ROW_43_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06653__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ net1344 net837 net816 _03354_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
XANTENNA__12217__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11240_ net882 net884 _05099_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11171_ net1341 net532 net525 _05073_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10122_ net1496 net172 net461 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XANTENNA__13037__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09355__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ net184 net2236 net424 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07905__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13812_ clknet_leaf_70_clk _01353_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10955_ net844 _04977_ top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__o21a_1
X_13743_ clknet_leaf_86_clk _01286_ net1016 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08330__B1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ clknet_leaf_103_clk _01232_ net1002 vssd1 vssd1 vccd1 vccd1 top.pc\[0\] sky130_fd_sc_hd__dfrtp_1
X_10886_ net1519 net228 net346 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
XANTENNA__07684__A2 _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06892__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ clknet_leaf_3_clk _00189_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ clknet_leaf_69_clk _00120_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06644__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ top.a1.dataIn\[15\] _05349_ _05371_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12487_ clknet_leaf_99_clk _00054_ net981 vssd1 vssd1 vccd1 vccd1 top.ramstore\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold109 net83 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _05301_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12424__Q top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10870__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _05223_ _05224_ _05212_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_210_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ clknet_leaf_45_clk _00672_ net1080 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13039_ clknet_leaf_21_clk _00603_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_206_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07600_ top.DUT.register\[6\]\[3\] net763 _02720_ _02726_ vssd1 vssd1 vccd1 vccd1
+ _02727_ sky130_fd_sc_hd__a211o_1
X_08580_ net270 _03494_ _03499_ net275 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_105_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07531_ top.DUT.register\[20\]\[4\] net578 net617 top.DUT.register\[30\]\[4\] _02648_
+ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ _02587_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__nand2_2
XANTENNA__10110__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07675__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ _04246_ _04247_ _04245_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06413_ net792 _01503_ _01506_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__and3_2
XANTENNA__06883__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07393_ _02186_ _02517_ _02206_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
X_09132_ _02690_ _02731_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__nand2_1
X_06344_ top.a1.instruction\[6\] _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07427__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06383__X _01510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06824__A _01929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06635__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _01992_ _02036_ _02077_ _02120_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__and4_1
X_06275_ top.ramload\[19\] net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[19\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__X _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ _03133_ _03135_ _03136_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__or4_1
Xhold610 top.DUT.register\[20\]\[5\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 top.DUT.register\[26\]\[22\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_116_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08388__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 top.DUT.register\[17\]\[5\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 top.DUT.register\[24\]\[25\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold654 top.DUT.register\[14\]\[5\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10780__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 top.DUT.register\[10\]\[10\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top.DUT.register\[4\]\[29\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 top.DUT.register\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07655__A _02759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 top.DUT.register\[11\]\[22\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net1369 net257 net429 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout582_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__C1 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ _03974_ _03994_ _04011_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__and3_1
X_09896_ net159 top.DUT.register\[1\]\[28\] net440 vssd1 vssd1 vccd1 vccd1 _00150_
+ sky130_fd_sc_hd__mux2_1
X_08847_ _03903_ _03946_ net281 vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__Y _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08778_ net521 _03879_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21ai_4
XANTENNA__13810__RESET_B net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07390__A top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ net287 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10020__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ net263 net1432 net375 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__mux2_1
XANTENNA__07666__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06874__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ net2223 net157 net452 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12410_ clknet_leaf_81_clk _00046_ net1006 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08933__B _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07418__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ clknet_leaf_117_clk _00954_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06734__A _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06626__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ _06132_ _06133_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12763__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12272_ _06091_ net1107 _06090_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__and3b_1
XFILLER_0_120_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11223_ net892 _05102_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__nor2_2
XANTENNA__10690__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09040__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ top.a1.state\[1\] net893 _04977_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_56_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11087__A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ net1521 net241 net459 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
X_11085_ net62 net859 vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_147_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08948__X _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ net246 net1711 net421 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__mux2_1
XANTENNA__11815__A top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08396__A _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06909__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11987_ _05799_ _05850_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ clknet_leaf_72_clk _01269_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_193_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10938_ net912 _04628_ _01416_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__or3b_2
XANTENNA__08854__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12419__Q top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10865__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ net464 _04942_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__nor2_8
X_13657_ clknet_leaf_91_clk _01216_ net998 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08606__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ clknet_leaf_46_clk _00172_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07409__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08606__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ clknet_leaf_97_clk _01147_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09020__A _03480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06617__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12539_ clknet_leaf_93_clk _00103_ net999 vssd1 vssd1 vccd1 vccd1 top.pc\[22\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07290__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12433__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07042__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 _04935_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_4
Xfanout419 _04927_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_6
XANTENNA__07593__A1 top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__B1 _03878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06962_ _02084_ _02086_ _02088_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__or3_1
XANTENNA__09961__Y _04920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ net833 _04356_ _04720_ top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _04758_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10105__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ _02950_ net468 net488 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__o21a_1
X_09681_ net835 _04199_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_1
X_06893_ top.DUT.register\[4\]\[22\] net565 net638 top.DUT.register\[16\]\[22\] _02019_
+ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a221o_1
XANTENNA__07481__Y _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _03076_ net487 net468 _03077_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__o22a_1
XANTENNA__07896__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ net284 _03468_ _03545_ _03409_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout163_A _04879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07514_ _01616_ _02639_ _02640_ net528 top.a1.instruction\[25\] vssd1 vssd1 vccd1
+ vccd1 _02641_ sky130_fd_sc_hd__a32o_4
XFILLER_0_159_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09689__X _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07648__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ _03555_ _03610_ _02448_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ top.DUT.register\[9\]\[6\] net629 net613 top.DUT.register\[14\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XANTENNA__06856__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10775__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout330_A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07376_ top.DUT.register\[6\]\[7\] net763 net693 top.DUT.register\[21\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _04172_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__nor2_1
X_06327_ _01457_ _01463_ _01335_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09046_ _03204_ _03295_ _03372_ net311 net319 vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o311a_1
XANTENNA__07281__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06258_ net1890 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[2\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout797_A _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold440 top.DUT.register\[20\]\[10\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07656__Y _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09022__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06189_ top.a1.halfData\[5\] _01416_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold451 top.DUT.register\[30\]\[12\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 top.DUT.register\[29\]\[19\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07033__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold473 top.DUT.register\[29\]\[22\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 top.DUT.register\[31\]\[24\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 top.DUT.register\[26\]\[27\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net934 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_2
Xfanout931 net933 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10015__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ net192 net1923 net436 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__mux2_1
Xfanout942 net946 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_2
Xfanout964 net980 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_2
Xfanout975 net977 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_4
Xfanout986 net996 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 net1020 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__buf_4
XANTENNA__13309__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _04869_ _04873_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_129_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 top.DUT.register\[5\]\[7\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 top.pad.keyCode\[4\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _05721_ _05764_ _05749_ net129 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a2bb2o_1
Xhold1162 top.DUT.register\[20\]\[17\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1173 top.DUT.register\[10\]\[2\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07887__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12890_ clknet_leaf_54_clk _00454_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_187_Left_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1184 top.DUT.register\[2\]\[29\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11841_ _05707_ _05710_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_142_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06448__B top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11772_ top.a1.dataIn\[8\] _05638_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07639__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06847__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ clknet_leaf_7_clk _01075_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10723_ net229 net1548 net384 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XANTENNA__09015__C_N _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10685__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10654_ net1704 net221 net452 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__mux2_1
X_13442_ clknet_leaf_49_clk _01006_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06464__A top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13373_ clknet_leaf_107_clk _00937_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10585_ net243 net1945 net387 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06183__B top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload18 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_4
Xclkload29 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload29/X sky130_fd_sc_hd__clkbuf_8
X_12324_ top.pad.button_control.debounce top.pad.button_control.noisy vssd1 vssd1
+ vccd1 vccd1 _06122_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07272__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07811__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12255_ top.lcd.cnt_20ms\[7\] top.lcd.cnt_20ms\[6\] _06065_ vssd1 vssd1 vccd1 vccd1
+ _06081_ sky130_fd_sc_hd__and3_1
XANTENNA__07024__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11206_ net850 _05076_ net531 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12186_ _06054_ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__or2_1
XANTENNA_hold4_A top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11137_ net60 net857 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07582__X _02709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ net1269 net862 net826 top.ramstore\[19\] vssd1 vssd1 vccd1 vccd1 _01186_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08524__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net185 net1654 net427 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
XANTENNA__07878__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__A _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07461__C _02586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06550__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06838__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ clknet_leaf_75_clk _01257_ net1091 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10595__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07230_ _02341_ _02352_ _02354_ _02356_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__nor4_1
XFILLER_0_184_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07161_ top.DUT.register\[28\]\[13\] net586 _01535_ top.DUT.register\[3\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07263__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ top.DUT.register\[23\]\[10\] net561 net600 top.DUT.register\[10\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12203__A2_N _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06369__A2 top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout216 net218 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlymetal6s2s_1
X_09802_ top.pc\[20\] _04443_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__or2_1
Xfanout227 net230 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
Xfanout238 _04723_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout249 _04707_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_1
X_07994_ top.DUT.register\[20\]\[31\] net749 net669 top.DUT.register\[5\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__a22o_1
X_06945_ top.DUT.register\[29\]\[21\] net665 net638 top.DUT.register\[16\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ net894 _04318_ _04741_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a21o_1
XANTENNA__09851__C _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ top.DUT.register\[9\]\[22\] net710 net677 top.DUT.register\[18\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
X_09664_ net465 _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__nand2_1
XANTENNA__07869__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08615_ net322 _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09595_ top.edg2.flip1 _01389_ _01604_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout545_A _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08546_ net479 _03656_ _03660_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06829__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08477_ net1303 net837 net818 _03594_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07428_ _02549_ _02551_ _02553_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__or4_2
XFILLER_0_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13398__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07359_ top.DUT.register\[20\]\[8\] net576 net603 top.DUT.register\[18\]\[8\] _02475_
+ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07254__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ net466 _04924_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ _04066_ _04090_ _03784_ _03896_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07006__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ top.a1.dataIn\[4\] _05877_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__nand2_1
Xhold270 top.DUT.register\[3\]\[16\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 top.DUT.register\[4\]\[31\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 top.a1.row2\[8\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout750 _01517_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_4
Xfanout761 _01510_ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout772 _01504_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_195_Left_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_4
Xfanout794 _01492_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_4
X_12942_ clknet_leaf_117_clk _00506_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ clknet_leaf_3_clk _00437_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08809__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11824_ _05679_ _05692_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__and2_1
XANTENNA__08674__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11755_ _05581_ _05615_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07493__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ net143 net1749 net379 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13425_ clknet_leaf_118_clk _00989_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09001__C net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10637_ net167 net2078 net392 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
Xclkload107 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__inv_4
XFILLER_0_141_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09709__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07245__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10568_ net189 net1615 net358 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__mux2_1
X_13356_ clknet_leaf_10_clk _00920_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ top.lcd.cnt_500hz\[10\] _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__or2_1
XANTENNA__07296__Y _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10499_ net213 top.DUT.register\[18\]\[18\] net368 vssd1 vssd1 vccd1 vccd1 _00684_
+ sky130_fd_sc_hd__mux2_1
X_13287_ clknet_leaf_7_clk _00851_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12238_ _06066_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__nor2_2
XANTENNA__12432__Q top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _06035_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
XANTENNA__07753__A _02879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06771__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06730_ top.DUT.register\[20\]\[26\] net579 net637 top.DUT.register\[16\]\[26\] _01844_
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a221o_1
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06661_ top.DUT.register\[8\]\[27\] net739 net731 top.DUT.register\[19\]\[27\] _01787_
+ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__inv_2
X_09380_ net821 _02519_ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__o21a_2
X_06592_ top.DUT.register\[20\]\[29\] net578 net657 top.DUT.register\[1\]\[29\] _01718_
+ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a221o_1
X_08331_ _03223_ _03230_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08262_ net481 net275 _03386_ _03382_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11280__A1 top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08871__X _03970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07213_ top.DUT.register\[1\]\[15\] net655 net615 top.DUT.register\[30\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__a22o_1
X_08193_ net278 _03315_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07144_ _02262_ _02264_ _02266_ _02270_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__or4_1
XANTENNA__07236__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06391__X _01518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ _01595_ _02187_ _02193_ _02200_ _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _01775_ _03103_ _01736_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout662_A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09716_ _03616_ net341 net338 _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__o211a_2
X_06928_ _02039_ _02041_ _02053_ _02054_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__or4_1
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ top.pc\[1\] _02788_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or2_1
X_06859_ top.DUT.register\[31\]\[23\] net743 net727 top.DUT.register\[10\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ top.pc\[30\] _04587_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12536__RESET_B net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08529_ _02277_ _03642_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08267__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _01393_ _05378_ net250 vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__nand3_1
XFILLER_0_203_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06445__C top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11471_ _05281_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire458 _04936_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
XANTENNA__07227__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ net240 net1627 net324 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__mux2_1
X_13210_ clknet_leaf_16_clk _00774_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08975__B1 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ clknet_leaf_6_clk _00705_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10353_ net1375 net229 net396 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__mux2_1
XANTENNA__07557__B _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06461__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ clknet_leaf_121_clk _00636_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10284_ net1383 net179 net401 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12023_ _05891_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__and2_1
XANTENNA__07844__Y _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13413__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout580 _01513_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06753__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout591 _04042_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_6
XANTENNA__10203__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ clknet_leaf_103_clk _00489_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ clknet_leaf_13_clk _00420_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _05672_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__nand2_2
XFILLER_0_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12787_ clknet_leaf_4_clk _00351_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07466__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ _05512_ _05541_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11262__B2 top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12427__Q top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11669_ _05534_ _05537_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13408_ clknet_leaf_45_clk _00972_ net1080 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07218__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__B1 _03072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13339_ clknet_leaf_48_clk _00903_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06371__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07900_ top.DUT.register\[15\]\[17\] net779 _03015_ _03026_ vssd1 vssd1 vccd1 vccd1
+ _03027_ sky130_fd_sc_hd__a211o_1
XANTENNA_max_cap513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08880_ _01778_ _03959_ _01776_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_4_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07831_ top.DUT.register\[11\]\[18\] net758 net695 top.DUT.register\[21\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a22o_1
XANTENNA__06744__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ _02608_ _02632_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_108_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09501_ _04535_ _04536_ _04537_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__and3_1
XFILLER_0_196_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06713_ _01833_ _01839_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__nor2_8
X_07693_ _02815_ _02817_ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__or3_1
XFILLER_0_211_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06644_ top.DUT.register\[1\]\[28\] net657 net565 top.DUT.register\[4\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22o_1
X_09432_ _04472_ _04473_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06575_ top.DUT.register\[20\]\[29\] net749 net746 top.DUT.register\[31\]\[29\] _01701_
+ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a221o_1
X_09363_ _04393_ _04397_ _04395_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout243_A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07457__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08314_ net886 top.pc\[3\] net536 _03437_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a22o_1
XANTENNA__11253__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ top.pc\[13\] _04318_ _04337_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08245_ net302 _03369_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10783__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13835__RESET_B net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07209__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11005__A1 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _02380_ net297 vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__or2_1
XANTENNA__12202__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08957__B1 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ _02239_ _02248_ _02251_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__nor4_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__X _03072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ top.a1.instruction\[28\] _01621_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06983__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08489__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10971_ top.a1.data\[0\] _04994_ _04989_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
X_12710_ clknet_leaf_24_clk _00274_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07696__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13690_ clknet_leaf_75_clk _01238_ net1088 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07160__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12641_ clknet_leaf_27_clk _00205_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07448__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ clknet_leaf_77_clk _00136_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11523_ _05349_ _05371_ _05368_ _05366_ _05363_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10693__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06472__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11454_ _05281_ _05317_ _05318_ _05322_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10405_ net176 net2304 net327 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__mux2_1
X_11385_ top.a1.dataIn\[30\] _05194_ _05249_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13124_ clknet_leaf_39_clk _00688_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09783__A top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10336_ net466 _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__nor2_1
XANTENNA__06974__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _04685_ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__nand2b_4
X_13055_ clknet_leaf_112_clk _00619_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08970__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _05828_ _05875_ _05845_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a21boi_1
X_10198_ net143 net1834 net410 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06726__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10868__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07750__B _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ clknet_leaf_9_clk _00472_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08884__C1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888_ net1138 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__09023__A _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_196_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ clknet_leaf_27_clk _00403_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06360_ net905 _01488_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__or2_2
XFILLER_0_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06291_ top.lcd.cnt_500hz\[9\] top.lcd.cnt_500hz\[11\] top.lcd.cnt_500hz\[10\] vssd1
+ vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__and3_1
XANTENNA__07749__Y _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08030_ _01579_ _01580_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap511 _02117_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold803 top.DUT.register\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold814 top.DUT.register\[24\]\[9\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 top.DUT.register\[12\]\[18\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10108__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold836 top.DUT.register\[13\]\[4\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 top.DUT.register\[26\]\[23\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold858 top.DUT.register\[22\]\[4\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ net1491 net203 net432 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
Xhold869 top.DUT.register\[11\]\[4\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _04025_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nand2_2
XFILLER_0_209_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08863_ _01776_ net468 net487 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__o21a_1
XANTENNA__06717__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ top.DUT.register\[19\]\[19\] net634 _01682_ top.DUT.register\[15\]\[19\]
+ _02929_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__a221o_1
X_08794_ net471 _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10778__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ top.DUT.register\[20\]\[1\] net749 net714 top.DUT.register\[30\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09667__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07678__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07676_ top.DUT.register\[28\]\[0\] net651 _02790_ _02802_ vssd1 vssd1 vccd1 vccd1
+ _02803_ sky130_fd_sc_hd__a211o_1
XANTENNA__07142__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _04455_ _04457_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__xnor2_1
X_06627_ _01742_ _01743_ _01751_ _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__or4_4
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout625_A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _03054_ _04378_ _04380_ _04381_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09868__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06558_ top.DUT.register\[1\]\[30\] net656 net564 top.DUT.register\[4\]\[30\] _01684_
+ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06489_ _01564_ net528 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _02255_ _04318_ _04321_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ net887 top.pc\[1\] net536 _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__a22o_1
XANTENNA__07850__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08159_ net516 net297 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__nand2_1
XANTENNA__10018__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07602__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ top.a1.dataInTemp\[7\] top.a1.data\[7\] net799 vssd1 vssd1 vccd1 vccd1 _05073_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06956__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net2008 net175 net459 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XANTENNA__07394__Y _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ net187 net2028 net424 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__mux2_1
XANTENNA__06708__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07381__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ clknet_leaf_70_clk net1163 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.debounce_dly
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10688__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06738__Y _01865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07669__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13742_ clknet_leaf_86_clk _01285_ net1016 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10954_ top.a1.halfData\[0\] _01379_ _01417_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__mux2_1
XANTENNA__07133__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__B2 _02685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ clknet_leaf_67_clk _01231_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10885_ net1549 net181 net346 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ clknet_leaf_0_clk _00188_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ clknet_leaf_69_clk _00119_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11506_ _05349_ _05371_ top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07841__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ clknet_leaf_114_clk _00053_ net981 vssd1 vssd1 vccd1 vccd1 top.ramstore\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11437_ _05302_ _05304_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nor3_1
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07585__X _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12193__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ _05236_ _05237_ _05232_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_210_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_1_clk _00671_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ net1470 net228 net400 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
X_11299_ _05093_ _05096_ _05160_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12639__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ clknet_leaf_117_clk _00602_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06929__X _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07372__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09649__A1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10598__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07530_ _02650_ _02652_ _02653_ _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__or4_1
XANTENNA__07124__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07461_ _02555_ _02561_ _02586_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__or3_2
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06412_ net790 _01503_ _01508_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__and3_4
X_09200_ _04254_ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07392_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06343_ top.a1.instruction\[2\] top.a1.instruction\[3\] _01473_ vssd1 vssd1 vccd1
+ vccd1 _01475_ sky130_fd_sc_hd__or3_2
X_09131_ _02690_ _02731_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09062_ _02448_ _02877_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nand2_1
XANTENNA__07832__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06274_ top.ramload\[18\] net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[18\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__13080__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08013_ top.DUT.register\[29\]\[31\] net665 net569 top.DUT.register\[8\]\[31\] _03139_
+ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold600 top.DUT.register\[25\]\[22\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold611 top.DUT.register\[26\]\[9\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout206_A _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold622 top.DUT.register\[9\]\[2\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__B2 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold633 top.DUT.register\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 top.DUT.register\[24\]\[0\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold655 top.DUT.register\[31\]\[6\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06399__B1 _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 top.DUT.register\[18\]\[2\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 top.DUT.register\[11\]\[2\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold688 top.DUT.register\[27\]\[13\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ net1382 net261 net429 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
Xhold699 top.DUT.register\[4\]\[0\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07655__B net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08915_ _03974_ _03994_ _04011_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a21oi_1
X_09895_ net337 _04880_ _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout575_A _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08846_ _01840_ net297 _03283_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07899__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08777_ net474 _03867_ _03870_ net471 _03880_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout742_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _02835_ _02854_ net806 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
XANTENNA__08312__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07115__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08312__B2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ _02785_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10670_ net1577 net161 net453 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09329_ _04373_ _04376_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07389__Y _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09273__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06734__B _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ net1855 _06130_ net795 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12271_ top.lcd.cnt_20ms\[13\] top.lcd.cnt_20ms\[12\] _06087_ vssd1 vssd1 vccd1 vccd1
+ _06091_ sky130_fd_sc_hd__and3_1
X_11222_ net883 _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09040__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ top.a1.row1\[101\] _04636_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__or2_1
XANTENNA__07565__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ net1636 net243 net460 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XANTENNA__11087__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ net915 net1344 net853 _05028_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ net252 net2270 net424 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XANTENNA__07354__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06909__B _02034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10211__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11986_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__inv_2
XANTENNA__09350__A_N _03012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ clknet_leaf_74_clk _01268_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfxtp_1
X_10937_ _00017_ _01416_ _04629_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_193_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08955__A1_N net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13656_ clknet_leaf_88_clk _01215_ net1006 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868_ net1461 net141 net351 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ clknet_leaf_113_clk _00171_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ clknet_leaf_98_clk _01146_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10799_ net1896 net158 net448 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09020__B _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ clknet_leaf_93_clk _00102_ net999 vssd1 vssd1 vccd1 vccd1 top.pc\[21\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07814__B1 _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10881__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12469_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[21\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[21\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07756__A _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout409 net412 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07593__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__B2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ top.DUT.register\[6\]\[20\] net766 net583 top.DUT.register\[12\]\[20\] _02087_
+ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ _02950_ net486 vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nand2_1
X_09680_ _04699_ top.DUT.register\[1\]\[3\] net437 vssd1 vssd1 vccd1 vccd1 _00125_
+ sky130_fd_sc_hd__mux2_1
X_06892_ top.DUT.register\[25\]\[22\] net626 net606 top.DUT.register\[18\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
X_08631_ net490 net521 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or2_2
XANTENNA__06553__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ net320 _03675_ _03674_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__o21a_1
XANTENNA__10121__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07513_ _02206_ _02609_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__or2_1
X_08493_ net503 _02447_ _02493_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout156_A _04890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07444_ top.DUT.register\[13\]\[6\] net650 net550 top.DUT.register\[24\]\[6\] _02568_
+ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a221o_1
XFILLER_0_186_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06394__X _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07375_ top.DUT.register\[19\]\[7\] net731 net704 top.DUT.register\[15\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout323_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ _04049_ _04175_ _04167_ _04166_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__a211o_1
X_06326_ _01450_ _01461_ _01466_ _01449_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07805__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10791__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ _03350_ _03389_ _03432_ _03446_ net319 vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o41a_1
X_06257_ net2102 net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[1\] sky130_fd_sc_hd__and2_1
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06188_ top.a1.halfData\[5\] _01416_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__or2_1
Xhold430 top.DUT.register\[18\]\[19\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09022__A2 _03426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold441 top.DUT.register\[7\]\[14\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 top.DUT.register\[11\]\[5\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 top.DUT.register\[11\]\[24\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 top.DUT.register\[22\]\[3\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 top.DUT.register\[10\]\[16\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 top.DUT.register\[29\]\[26\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 net911 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_2
Xfanout921 net934 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
X_09947_ net204 net2081 net436 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__mux2_1
Xfanout943 net946 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_2
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
XANTENNA_fanout957_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net968 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
Xfanout976 net977 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
Xfanout987 net989 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_4
X_09878_ _04869_ _04873_ net804 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_129_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 top.DUT.register\[10\]\[13\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
Xhold1141 top.DUT.register\[30\]\[22\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07336__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__A3 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ net300 _03929_ _03927_ net269 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__o211a_1
Xhold1152 top.DUT.register\[4\]\[8\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 top.DUT.register\[5\]\[18\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 top.DUT.register\[21\]\[29\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ _05673_ _05708_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10031__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11771_ _05603_ _05637_ _05639_ _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_178_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08836__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ clknet_leaf_20_clk _01074_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10722_ net182 net1394 net381 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09121__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ clknet_leaf_25_clk _01005_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ net1416 net226 net453 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13372_ clknet_leaf_54_clk _00936_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10584_ net247 net2175 net386 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
Xclkload19 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ net912 net118 _06120_ top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 _01352_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07272__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09549__B1 _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ top.lcd.cnt_20ms\[6\] _06065_ top.lcd.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ _06080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ net1209 net530 _05089_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_71_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10206__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12185_ top.a1.dataIn\[1\] _06050_ _06052_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__and3_1
XANTENNA__07575__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__X _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ net917 net2141 net852 _05054_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a31o_1
XANTENNA__06783__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11067_ net82 net862 net827 net1239 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07327__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12694__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ net189 net2010 net427 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XANTENNA__09015__B _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10876__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11969_ _05811_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__xnor2_2
X_13708_ clknet_leaf_73_clk _01256_ net1093 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12541__SET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13639_ clknet_leaf_45_clk net1234 net1081 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07160_ top.DUT.register\[4\]\[13\] net768 net715 top.DUT.register\[30\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08202__A1_N net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ top.DUT.register\[17\]\[10\] net643 net619 top.DUT.register\[26\]\[10\] _02217_
+ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10116__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 _04802_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
X_09801_ top.pc\[20\] _04443_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__and2_1
XANTENNA__07566__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 net230 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkload10_A clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout239 net242 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
X_07993_ top.DUT.register\[4\]\[31\] net769 _03114_ _03119_ vssd1 vssd1 vccd1 vccd1
+ _03120_ sky130_fd_sc_hd__a211o_1
XANTENNA__06774__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ net894 _04318_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__and3_1
X_06944_ top.DUT.register\[21\]\[21\] net574 net553 top.DUT.register\[7\]\[21\] _02070_
+ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a221o_1
XANTENNA__06389__X _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11114__A3 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09712__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _04678_ _04685_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nor2_1
XANTENNA__08110__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ top.DUT.register\[27\]\[22\] net778 net766 top.DUT.register\[6\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout273_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _03538_ _03725_ net310 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09594_ net908 top.pc\[31\] _04618_ _04626_ net897 vssd1 vssd1 vccd1 vccd1 _00112_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_210_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08545_ _02275_ net486 net478 _03658_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout440_A _04681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ net887 top.pc\[9\] net536 _03593_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a22o_1
XANTENNA__06565__A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07427_ top.DUT.register\[20\]\[6\] net750 net725 top.DUT.register\[17\]\[6\] _02546_
+ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout705_A _01533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07358_ _02477_ _02479_ _02480_ _02484_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06309_ _01452_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07289_ top.DUT.register\[22\]\[9\] net752 net705 top.DUT.register\[15\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09028_ _03619_ _03830_ _04089_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 top.DUT.register\[19\]\[23\] vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 top.DUT.register\[29\]\[29\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 top.DUT.register\[26\]\[13\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 top.ramaddr\[26\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06765__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 _01519_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_2
Xfanout751 _01516_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_8
Xfanout762 _01510_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07309__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout784 _01659_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
Xfanout795 _06124_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09116__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ clknet_leaf_25_clk _00505_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__B net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ clknet_leaf_35_clk _00436_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07190__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08809__A2 _03742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11754_ _05574_ _05622_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06475__A _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10268__Y _04939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10705_ net146 net2105 net378 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ _05522_ _05553_ _05519_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13424_ clknet_leaf_2_clk _00988_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ net168 net1995 net390 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13355_ clknet_leaf_31_clk _00919_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10567_ net194 net2048 net359 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12306_ _06111_ net588 _06110_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__and3b_1
XANTENNA__07796__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ clknet_leaf_19_clk _00850_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_188_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10498_ net216 net2208 net365 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _06067_ _06068_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__or3_1
XANTENNA__07548__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ _06027_ net125 _06033_ _06036_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o22ai_1
XANTENNA__06756__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11119_ net50 net859 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_207_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12099_ _05968_ _05940_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__and2b_1
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06660_ top.DUT.register\[27\]\[27\] net775 net697 top.DUT.register\[23\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07181__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_max_cap493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__C1 top.i_ready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06591_ top.DUT.register\[24\]\[29\] net550 net617 top.DUT.register\[30\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08330_ _02684_ _03177_ net469 _02685_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_59_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08076__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08261_ net304 _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__nand2_2
XFILLER_0_46_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07212_ _02331_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__nor2_4
XANTENNA_wire496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08804__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08192_ net278 _03316_ _03317_ net300 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07143_ top.DUT.register\[23\]\[12\] net563 net558 top.DUT.register\[6\]\[12\] _02269_
+ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08433__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _01481_ _01576_ _01478_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1028_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout390_A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _01778_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__or2_1
X_09715_ top.pc\[10\] net803 _04718_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a211o_1
X_06927_ top.DUT.register\[6\]\[21\] net766 net682 top.DUT.register\[7\]\[21\] _02051_
+ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout655_A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ top.a1.halfData\[5\] _01472_ _04658_ net1105 vssd1 vssd1 vccd1 vccd1 _00120_
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_27_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06858_ top.DUT.register\[29\]\[23\] net700 _01954_ _01984_ vssd1 vssd1 vccd1 vccd1
+ _01985_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07172__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07711__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_182_Right_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09577_ _04598_ _04599_ _04596_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_26_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ top.DUT.register\[6\]\[24\] net765 net698 top.DUT.register\[23\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08528_ _02277_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06445__D top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11470_ _05308_ _05319_ _05321_ net267 _05311_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a41o_1
XANTENNA_clkbuf_4_6__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10421_ net245 top.DUT.register\[16\]\[6\] net326 vssd1 vssd1 vccd1 vccd1 _00608_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ clknet_leaf_47_clk _00704_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08975__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10352_ net1545 net181 net393 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13071_ clknet_leaf_20_clk _00635_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ net1502 net196 net403 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12022_ _05868_ net127 _05871_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_4
Xfanout581 _01513_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_2
Xfanout592 _04042_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_45_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12924_ clknet_leaf_53_clk _00488_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07163__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ clknet_leaf_107_clk _00419_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12202__A2_N _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _05662_ _05673_ _05675_ _05674_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__o31a_2
XFILLER_0_56_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12786_ clknet_leaf_52_clk _00350_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08570__A2_N net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11737_ _05547_ _05567_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11668_ _05534_ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_54_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13407_ clknet_leaf_113_clk _00971_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ net236 net2226 net389 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__mux2_1
XANTENNA__12211__A1 top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11599_ _05457_ _05462_ _05465_ _05466_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13338_ clknet_leaf_15_clk _00902_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08966__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06977__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13269_ clknet_leaf_6_clk _00833_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08212__X _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07830_ top.DUT.register\[27\]\[18\] net778 net738 top.DUT.register\[24\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07761_ _02636_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__nand2_1
X_09500_ _04536_ _04537_ _04535_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a21oi_1
X_06712_ _01827_ _01828_ _01836_ _01838_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_108_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07692_ top.DUT.register\[19\]\[0\] net731 net704 top.DUT.register\[15\]\[0\] _02818_
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a221o_1
XANTENNA__07154__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ top.pc\[22\] _04460_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06643_ top.DUT.register\[24\]\[28\] net551 net542 top.DUT.register\[22\]\[28\] _01769_
+ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a221o_1
XANTENNA__06386__Y _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ _02970_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09203__B _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06574_ top.DUT.register\[27\]\[29\] net777 net729 top.DUT.register\[10\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ _03434_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__nand2_2
X_09293_ _04341_ _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_72_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ _03193_ _03200_ net287 vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11005__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08175_ _02298_ net297 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nand2_1
XANTENNA__06680__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout403_A _04939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08957__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07126_ top.DUT.register\[11\]\[12\] net757 net706 top.DUT.register\[15\]\[12\] _02252_
+ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a221o_1
XANTENNA__06968__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07057_ _02175_ _02183_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__nor2_8
XFILLER_0_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10304__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _02951_ _03085_ _03080_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ top.a1.dataIn\[0\] net849 _04990_ _04993_ vssd1 vssd1 vccd1 vccd1 _04994_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07145__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _04645_ _04651_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__nor2_1
XANTENNA__06499__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06296__Y _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ clknet_leaf_49_clk _00204_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08645__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ clknet_leaf_56_clk _00135_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_50_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11522_ _05365_ _05391_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11453_ _05281_ _05318_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__nor3_1
XANTENNA__06671__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ net183 net2178 net329 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11384_ _05251_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__and2b_1
XANTENNA__06959__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13123_ clknet_leaf_22_clk _00687_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10335_ _04916_ _04937_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09783__B _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06423__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ clknet_leaf_13_clk _00618_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ top.a1.instruction\[9\] top.a1.instruction\[10\] _04675_ vssd1 vssd1 vccd1
+ vccd1 _04937_ sky130_fd_sc_hd__and3_2
X_12005_ _05840_ _05844_ _05825_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a21o_1
XANTENNA__10214__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10197_ net145 net1540 net412 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07384__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07923__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07136__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12907_ clknet_leaf_30_clk _00471_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13887_ net1137 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10691__A0 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09798__X _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12838_ clknet_leaf_20_clk _00402_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_196_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07439__A1 top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ clknet_leaf_28_clk _00333_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06290_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[3\] top.lcd.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06662__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12196__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold804 top.DUT.register\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 top.DUT.register\[12\]\[13\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold826 top.DUT.register\[23\]\[6\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold837 top.DUT.register\[25\]\[24\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 top.DUT.register\[7\]\[23\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ net2268 net211 net431 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
Xhold859 top.DUT.register\[26\]\[31\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ net475 _04017_ _04018_ net472 _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__o221a_1
XFILLER_0_149_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13215__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ _03191_ _03199_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nand2_1
XANTENNA__10124__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07914__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ top.DUT.register\[20\]\[19\] net578 net628 top.DUT.register\[9\]\[19\] _02939_
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a221o_1
X_08793_ _01953_ _03095_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout186_A _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07744_ top.DUT.register\[23\]\[1\] net698 net672 top.DUT.register\[16\]\[1\] _02870_
+ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a221o_1
XANTENNA__09667__A2 _01492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07675_ top.DUT.register\[19\]\[0\] net631 net781 top.DUT.register\[31\]\[0\] _02801_
+ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout353_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12850__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ _04439_ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1095_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06626_ top.DUT.register\[17\]\[28\] net724 net717 top.DUT.register\[2\]\[28\] _01752_
+ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__a221o_1
XFILLER_0_181_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _04390_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout520_A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06557_ top.DUT.register\[29\]\[30\] net664 net781 top.DUT.register\[31\]\[30\] _01683_
+ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout618_A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08772__B net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06488_ net833 net534 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__or2_4
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08227_ _03346_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06653__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07109_ _02165_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__nand2_1
X_08089_ net290 _03012_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10120_ net1895 net183 net460 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09355__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ net194 net1743 net423 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__mux2_1
XANTENNA__10034__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09346__A1_N _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07905__A2 _03031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ clknet_leaf_70_clk _00017_ net1106 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.noisy
+ sky130_fd_sc_hd__dfrtp_1
X_13889__1139 vssd1 vssd1 vccd1 vccd1 _13889__1139/HI net1139 sky130_fd_sc_hd__conb_1
XANTENNA__07118__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ clknet_leaf_86_clk _01284_ net1016 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_119_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10953_ _01410_ _04979_ _04982_ _04981_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13642__Q net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06467__B top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ clknet_leaf_95_clk net1164 net988 vssd1 vssd1 vccd1 vccd1 wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ net2165 net198 net347 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12520__RESET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12623_ clknet_leaf_20_clk _00187_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06892__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ clknet_leaf_69_clk _00118_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _05337_ _05372_ _05373_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06644__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12485_ clknet_leaf_61_clk _00052_ net1099 vssd1 vssd1 vccd1 vccd1 top.ramstore\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10209__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11436_ _05263_ _05292_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_128_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11232__A_N net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11367_ _05207_ _05233_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__xor2_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ clknet_leaf_51_clk _00670_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ net2194 net181 net397 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
X_11298_ net1194 net824 _05172_ net1093 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_165_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ clknet_leaf_23_clk _00601_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ net1372 net180 net455 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__mux2_1
XANTENNA__10879__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08857__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07460_ _02562_ _02586_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06411_ top.DUT.register\[11\]\[30\] net756 net697 top.DUT.register\[23\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06883__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ top.a1.instruction\[19\] _01617_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08592__B _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ _04187_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__xnor2_1
X_06342_ top.a1.instruction\[3\] _01473_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09061_ _03378_ _03514_ _03610_ _03662_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__and4_1
XANTENNA__06635__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06273_ top.ramload\[17\] net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[17\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_72_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10119__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13467__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08012_ top.DUT.register\[15\]\[31\] _01682_ _03137_ _03138_ vssd1 vssd1 vccd1 vccd1
+ _03139_ sky130_fd_sc_hd__a211o_1
Xhold601 top.DUT.register\[16\]\[23\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 top.DUT.register\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap331 _05283_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_116_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 top.DUT.register\[23\]\[2\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 top.DUT.register\[8\]\[29\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 top.DUT.register\[31\]\[23\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 top.DUT.register\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07596__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 top.DUT.register\[15\]\[13\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 top.DUT.register\[18\]\[3\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net1487 net263 net432 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__mux2_1
XANTENNA__08113__A _02339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 top.DUT.register\[5\]\[14\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09337__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _01692_ net485 _04010_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__a21boi_1
X_09894_ _04885_ _04886_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a21o_1
XANTENNA__07348__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08845_ net309 _03873_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__or2_1
XANTENNA__10789__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout470_A _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _03533_ _03771_ _03875_ net482 _03877_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__o221a_1
XFILLER_0_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07727_ _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_A _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07658_ net902 net524 _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07520__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06609_ _01734_ _01735_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06874__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_A top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ top.DUT.register\[25\]\[3\] net772 net747 top.DUT.register\[20\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09328_ _04374_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06626__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09259_ net911 top.pc\[11\] _04311_ net899 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12270_ top.lcd.cnt_20ms\[12\] top.lcd.cnt_20ms\[11\] _06086_ top.lcd.cnt_20ms\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ net879 top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07587__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _01432_ _01435_ _05063_ top.busy_o vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__o22a_1
XANTENNA__07051__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ net1709 net246 net459 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XANTENNA__12541__Q top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083_ net51 net859 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__and2_1
XANTENNA__07339__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10034_ net257 net1949 net421 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__mux2_1
XANTENNA__10699__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__Y _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12701__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11985_ _05844_ _05853_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10936_ top.a1.halfData\[5\] _01424_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__nand2_1
X_13724_ clknet_leaf_73_clk _01267_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13655_ clknet_leaf_87_clk _01214_ net1008 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
X_10867_ net1517 net144 net350 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ clknet_leaf_12_clk _00170_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13586_ clknet_leaf_95_clk _01145_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ net1660 net161 net446 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06617__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ clknet_leaf_90_clk _00101_ net999 vssd1 vssd1 vccd1 vccd1 top.pc\[20\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09728__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12468_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[20\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[20\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07290__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11419_ _05273_ _05283_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__a211o_2
XANTENNA__09567__B2 _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12399_ clknet_leaf_90_clk _00035_ net998 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07042__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09319__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09319__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ top.DUT.register\[29\]\[20\] net703 net694 top.DUT.register\[21\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_3_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11126__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06891_ top.DUT.register\[15\]\[22\] _01655_ net783 top.DUT.register\[31\]\[22\]
+ _02017_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a221o_1
X_08630_ net322 _03221_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10402__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ net284 _03483_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07512_ _02207_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__or2_1
X_08492_ _03183_ _03606_ _03608_ net480 vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07443_ top.DUT.register\[15\]\[6\] _01655_ net783 top.DUT.register\[31\]\[6\] _02569_
+ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06856__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout149_A _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ top.DUT.register\[3\]\[7\] net689 net684 top.DUT.register\[7\]\[7\] _02500_
+ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _04173_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__nand2_1
X_06325_ _01462_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11062__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1058_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09044_ _03484_ _03511_ _03533_ net314 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__a31o_1
X_06256_ net1340 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[0\] sky130_fd_sc_hd__and2_1
XANTENNA__07281__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888__1138 vssd1 vssd1 vccd1 vccd1 _13888__1138/HI net1138 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_131_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold420 top.DUT.register\[6\]\[7\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ _01413_ _01414_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__and2_1
Xhold431 top.DUT.register\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07569__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 top.pc\[0\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold453 top.DUT.register\[17\]\[10\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold464 top.DUT.register\[29\]\[8\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 top.ramload\[22\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 top.DUT.register\[21\]\[11\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__buf_2
XANTENNA_fanout685_A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout911 top.i_ready vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
Xhold497 top.DUT.register\[21\]\[4\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_4
X_09946_ net211 net1847 net436 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__mux2_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net946 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net980 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07682__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout966 net968 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08130__X _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _04870_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__nand2_1
Xhold1120 top.DUT.register\[5\]\[10\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 top.DUT.register\[7\]\[0\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
Xhold1142 top.a1.row2\[16\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _03888_ _03928_ net277 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__mux2_1
XANTENNA__10312__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1153 top.DUT.register\[2\]\[31\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 top.DUT.register\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06298__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12496__CLK clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07741__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1175 top.DUT.register\[10\]\[19\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 top.DUT.register\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ net475 _03851_ _03863_ net471 _03862_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__o221ai_4
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _05560_ _05620_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__or2_1
X_10721_ net198 net1552 net384 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06847__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13440_ clknet_leaf_45_clk _01004_ net1082 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_175_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10652_ net1498 net233 net451 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12536__Q top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13371_ clknet_leaf_52_clk _00935_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10583_ net252 net1657 net387 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ _06120_ _06121_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07272__A2 _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12253_ _01382_ _06066_ _06079_ net1108 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ net850 _05075_ net531 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__and3_1
XANTENNA__07024__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12184_ _06050_ _06052_ top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_71_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12953__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ net59 net857 vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_196_Right_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11066_ net1260 net856 net825 top.ramstore\[17\] vssd1 vssd1 vccd1 vccd1 _01184_
+ sky130_fd_sc_hd__a22o_1
X_10017_ net193 net2308 net427 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10222__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12989__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06495__X _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _05822_ _05823_ _05802_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13707_ clknet_leaf_73_clk _01255_ net1094 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06838__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ net227 net1477 net442 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
X_11899_ top.a1.dataIn\[5\] _05684_ _05729_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__or3_1
XANTENNA__09031__B _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13638_ clknet_leaf_45_clk net1310 net1081 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12446__Q top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10892__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13569_ clknet_leaf_84_clk _01128_ net1017 vssd1 vssd1 vccd1 vccd1 top.a1.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07090_ top.DUT.register\[11\]\[10\] net639 net607 top.DUT.register\[12\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
XANTENNA__07263__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08869__Y _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ top.pc\[19\] _04425_ _04797_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a21o_1
Xfanout207 net210 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
Xfanout218 _04786_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
Xfanout229 net230 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
X_07992_ top.DUT.register\[28\]\[31\] net586 net722 top.DUT.register\[14\]\[31\] _03118_
+ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09731_ _04739_ _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__nor2_1
X_06943_ top.DUT.register\[8\]\[21\] net570 net546 top.DUT.register\[5\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09712__A1 _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ top.a1.instruction\[7\] top.a1.instruction\[8\] _04675_ vssd1 vssd1 vccd1
+ vccd1 _04685_ sky130_fd_sc_hd__o21a_1
X_06874_ top.DUT.register\[28\]\[22\] net587 _01535_ top.DUT.register\[3\]\[22\] _02000_
+ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a221o_1
XANTENNA__08110__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _03622_ _03724_ net307 vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__mux2_1
X_09593_ net133 _04622_ _04623_ net137 net909 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_179_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout266_A _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ _02277_ net470 _03652_ net522 _03653_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_210_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06829__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ net472 _03575_ _03592_ net477 _03590_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_175_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout433_A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13740__Q top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07426_ top.DUT.register\[1\]\[6\] net688 net680 top.DUT.register\[13\]\[6\] _02552_
+ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07357_ top.DUT.register\[27\]\[8\] net595 _02482_ _02483_ vssd1 vssd1 vccd1 vccd1
+ _02484_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout600_A _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06308_ net1542 _01445_ _01446_ net883 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07254__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ top.DUT.register\[19\]\[9\] net732 net728 top.DUT.register\[10\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10374__Y _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06462__B1 _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09027_ _03645_ _03762_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nand2_1
XANTENNA__11199__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06239_ top.ramload\[15\] net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[15\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__13294__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07006__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 top.DUT.register\[28\]\[24\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold261 top.DUT.register\[7\]\[4\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 top.DUT.register\[26\]\[1\] vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 top.DUT.register\[28\]\[3\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top.DUT.register\[19\]\[20\] vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07683__Y _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout730 _01523_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 _01519_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_8
Xfanout752 _01516_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ net265 net2235 net435 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__mux2_1
Xfanout763 _01509_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 _01504_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
Xfanout785 _01657_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_4
XANTENNA__09703__A1 _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout796 _06124_ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10042__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12940_ clknet_leaf_8_clk _00504_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07714__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09831__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ clknet_leaf_7_clk _00435_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07190__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11822_ _05650_ _05690_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09132__A _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _05589_ _05600_ _05594_ _05574_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08019__Y _03146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10704_ net152 net2124 net379 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
X_11684_ _05519_ _05522_ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__and3_1
XANTENNA__07493__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ net171 net2265 net391 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__mux2_1
X_13423_ clknet_leaf_23_clk _00987_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13354_ clknet_leaf_38_clk _00918_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10566_ net203 net2287 net358 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__mux2_1
XANTENNA__07245__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ top.lcd.cnt_500hz\[9\] _06109_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__and2_1
X_13285_ clknet_leaf_120_clk _00849_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10217__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10497_ net227 net1677 net366 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ top.lcd.cnt_20ms\[15\] top.lcd.cnt_20ms\[14\] top.lcd.cnt_20ms\[17\] top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__or4bb_1
X_12167_ _06035_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11118_ net914 net1262 net853 _05045_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a31o_1
XANTENNA_output62_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872__1159 vssd1 vssd1 vccd1 vccd1 net1159 _13872__1159/LO sky130_fd_sc_hd__conb_1
X_12098_ _05956_ _05964_ _05955_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_207_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ net73 net860 net829 net1214 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a22o_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10887__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887__1137 vssd1 vssd1 vccd1 vccd1 _13887__1137/HI net1137 sky130_fd_sc_hd__conb_1
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06590_ top.DUT.register\[6\]\[29\] net558 net621 top.DUT.register\[26\]\[29\] _01716_
+ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ net287 _03384_ _03383_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07211_ _02333_ _02335_ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__or3_2
XFILLER_0_116_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08191_ net495 net289 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_99_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07142_ top.DUT.register\[15\]\[12\] net780 _02267_ _02268_ vssd1 vssd1 vccd1 vccd1
+ _02269_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07236__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__B2 _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07073_ _01571_ _01596_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__or2_1
XANTENNA__10127__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__Y _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07944__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__A _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _01797_ _01817_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06926_ top.DUT.register\[24\]\[21\] net738 net702 top.DUT.register\[29\]\[21\] _02052_
+ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a221o_1
X_09714_ net835 _04282_ _04720_ top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 _04727_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_126_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09697__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ _04667_ _04668_ _04669_ _04670_ net1106 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__o311a_1
XANTENNA__10797__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06857_ top.DUT.register\[21\]\[23\] net692 net681 top.DUT.register\[7\]\[23\] _01983_
+ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout550_A _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout648_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09576_ _01618_ _04608_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__and3_1
X_06788_ top.DUT.register\[31\]\[24\] net745 net741 top.DUT.register\[8\]\[24\] _01914_
+ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10369__Y _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11256__B1 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ _02906_ _03641_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__and2_1
XFILLER_0_194_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout815_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ _03280_ _03312_ net311 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07475__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07409_ top.DUT.register\[16\]\[7\] net636 net555 top.DUT.register\[7\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XANTENNA__11008__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06683__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08389_ _02589_ net469 _03508_ net481 _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ net247 net2057 net323 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__mux2_1
Xwire449 _04950_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_2
XFILLER_0_123_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08975__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ net1409 net198 net395 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__mux2_1
XANTENNA__10037__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13070_ clknet_leaf_111_clk _00634_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10282_ net1975 net200 net404 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12021_ _05868_ _05871_ _05878_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__nand3_1
XANTENNA__08302__Y _03426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13645__Q net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _01650_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09137__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout571 _01646_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_8
Xfanout582 _01513_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_8
Xfanout593 _04041_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_100_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12923_ clknet_leaf_48_clk _00487_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08360__B1 _03480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10500__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ clknet_leaf_119_clk _00418_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ _05613_ _05671_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12785_ clknet_leaf_116_clk _00349_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11736_ _05547_ _05572_ _05589_ _05599_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nor4_1
XANTENNA__07466__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08663__A1 _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06674__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ _05507_ _05535_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__xor2_1
XANTENNA__06492__Y _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ clknet_leaf_12_clk _00970_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07218__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10618_ net240 net1525 net390 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__mux2_1
XANTENNA__08206__A _02879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _05457_ _05462_ _05465_ _05466_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__and4bb_1
XANTENNA__12211__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08966__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13337_ clknet_leaf_36_clk _00901_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10549_ net259 net2317 net357 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13268_ clknet_leaf_46_clk _00832_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12219_ net1168 _06059_ net589 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
X_13199_ clknet_leaf_22_clk _00763_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09037__A _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire449_A _04950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07760_ net313 _02682_ _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09679__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ top.DUT.register\[28\]\[26\] net587 net702 top.DUT.register\[29\]\[26\] _01837_
+ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07691_ top.DUT.register\[26\]\[0\] net759 net712 top.DUT.register\[30\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09430_ top.pc\[22\] _04460_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nand2_1
X_06642_ top.DUT.register\[2\]\[28\] net661 net546 top.DUT.register\[5\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10410__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13074__RESET_B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ _01615_ _02519_ _02563_ net821 _01622_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__o221a_2
XTAP_TAPCELL_ROW_121_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06573_ top.DUT.register\[22\]\[29\] net753 _01535_ top.DUT.register\[3\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08312_ net519 _03412_ _03417_ net473 _03435_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07457__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ top.pc\[14\] _04325_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__nor2_1
X_08243_ net285 _03367_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__nor2_1
XANTENNA__06665__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout229_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08174_ net286 _03298_ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07209__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__A _02298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ top.DUT.register\[26\]\[12\] net761 net754 top.DUT.register\[22\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XANTENNA__08957__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _02176_ _02178_ _02180_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout598_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09367__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07917__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _02971_ _02990_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_199_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06909_ net514 _02034_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ top.DUT.register\[13\]\[17\] net647 net639 top.DUT.register\[11\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ top.a1.halfData\[0\] _01472_ _04656_ net1103 vssd1 vssd1 vccd1 vccd1 _00116_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10320__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06499__A3 _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _01619_ _04591_ _04592_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ clknet_leaf_15_clk _00134_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07448__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08645__B2 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09410__A top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ _05349_ _05371_ _05363_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_61_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06656__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871__1158 vssd1 vssd1 vccd1 vccd1 net1158 _13871__1158/LO sky130_fd_sc_hd__conb_1
XFILLER_0_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ _05280_ _05309_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_152_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08026__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10403_ net190 net2144 net330 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11383_ _05220_ _05224_ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13886__1136 vssd1 vssd1 vccd1 vccd1 _13886__1136/HI net1136 sky130_fd_sc_hd__conb_1
X_13122_ clknet_leaf_44_clk _00686_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10334_ net1882 net140 net398 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__mux2_1
XANTENNA__07865__A _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07620__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ clknet_leaf_108_clk _00617_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ net1581 net140 net456 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__mux2_1
X_12004_ _05860_ _05861_ _05864_ _05867_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a41oi_4
XTAP_TAPCELL_ROW_167_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10196_ net154 net1809 net410 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout390 _04944_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_4
XFILLER_0_108_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12906_ clknet_leaf_38_clk _00470_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10230__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ net1136 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_198_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06895__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_196_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12837_ clknet_leaf_118_clk _00401_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12768_ clknet_leaf_42_clk _00332_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06647__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__B _02685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ _05586_ _05588_ _05587_ _05563_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__o211a_2
XFILLER_0_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ clknet_leaf_47_clk _00263_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold805 top.DUT.register\[21\]\[22\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_2
XFILLER_0_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold816 top.DUT.register\[23\]\[7\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold827 top.DUT.register\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold838 top.DUT.register\[15\]\[0\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 top.DUT.register\[2\]\[11\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _03183_ _04023_ _03771_ _03719_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10405__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ _01778_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_209_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07812_ top.DUT.register\[2\]\[19\] net662 net625 top.DUT.register\[25\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a22o_1
X_08792_ _03892_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__or3b_2
XANTENNA__09054__X _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ top.DUT.register\[26\]\[1\] net761 net691 top.DUT.register\[3\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a22o_1
XANTENNA__08738__A1_N net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ top.DUT.register\[3\]\[0\] net785 net779 top.DUT.register\[15\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
XANTENNA__10140__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06625_ top.DUT.register\[6\]\[28\] net765 net758 top.DUT.register\[11\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
X_09413_ _04438_ _04440_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout346_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09344_ _04373_ _04374_ _04375_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__o21ai_1
X_06556_ top.DUT.register\[19\]\[30\] net632 net780 top.DUT.register\[15\]\[30\] _01658_
+ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_205_Left_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06638__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ net894 _04293_ top.pc\[13\] vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10376__A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06487_ net833 net534 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ net519 _03329_ _03351_ net479 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_43_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07850__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _01797_ net292 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10198__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07108_ _02233_ _02234_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__nand2_2
X_08088_ net295 _03054_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__nand2_1
XANTENNA__08133__X _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07602__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__A2_N _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ top.DUT.register\[8\]\[10\] net740 net668 top.DUT.register\[5\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XANTENNA__06810__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10315__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ net205 net2279 net423 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__C1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08315__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09512__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ clknet_leaf_85_clk _01283_ net1018 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10050__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ top.a1.hexop\[4\] _01417_ _01424_ _01384_ vssd1 vssd1 vccd1 vccd1 _04982_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07669__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12539__Q top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06877__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13671_ clknet_leaf_83_clk _01230_ net1017 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10883_ net2038 net201 net347 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12622_ clknet_leaf_111_clk _00186_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06629__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12553_ clknet_leaf_69_clk _00117_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08027__Y _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11504_ top.a1.dataIn\[15\] _05297_ _05334_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__or3_1
XANTENNA__07841__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12484_ clknet_leaf_83_clk _00051_ net1013 vssd1 vssd1 vccd1 vccd1 top.ramstore\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11435_ _05302_ _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07866__Y _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07054__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ top.a1.dataIn\[18\] _05233_ _05234_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_210_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13105_ clknet_leaf_3_clk _00669_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10317_ net1527 net195 net398 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__mux2_1
XANTENNA__10225__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ _05098_ _05171_ _05155_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__or3b_1
X_13036_ clknet_leaf_8_clk _00600_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10248_ net1489 net198 net455 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__mux2_1
XANTENNA__08554__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__C1 _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06498__X _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ net208 net1963 net410 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_198_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06580__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08857__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8__f_clk_X clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10895__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ net1156 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
X_06410_ _01497_ net792 _01506_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and3_4
XFILLER_0_201_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ top.a1.instruction\[27\] _01621_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06341_ top.a1.instruction\[0\] top.a1.instruction\[1\] vssd1 vssd1 vccd1 vccd1 _01473_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _04118_ _04119_ _04121_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__and3_1
X_06272_ top.ramload\[16\] net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[16\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07293__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ top.DUT.register\[28\]\[31\] net653 net634 top.DUT.register\[19\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a22o_1
Xhold602 top.DUT.register\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 top.DUT.register\[6\]\[25\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 top.DUT.register\[26\]\[28\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold635 top.DUT.register\[20\]\[13\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06399__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 top.DUT.register\[6\]\[30\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 top.DUT.register\[22\]\[5\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 top.DUT.register\[28\]\[26\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10135__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09962_ net1901 net151 net429 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
Xhold679 top.DUT.register\[26\]\[16\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09924__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ net475 _03998_ _03999_ net472 _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o221a_1
X_09893_ net835 _04568_ _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_209_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _03101_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__nand2_1
XANTENNA__07899__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870__1157 vssd1 vssd1 vccd1 vccd1 net1157 _13870__1157/LO sky130_fd_sc_hd__conb_1
X_08775_ net317 _03532_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__o21ba_2
XANTENNA__13743__Q top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout463_A _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07016__Y _02143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ _02848_ _02850_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nor3_1
XANTENNA__08848__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06859__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13885__1135 vssd1 vssd1 vccd1 vccd1 _13885__1135/HI net1135 sky130_fd_sc_hd__conb_1
X_07657_ top.a1.instruction\[8\] _01477_ _01620_ top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 _02784_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout728_A _01523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ _01713_ _01732_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__and2_1
XANTENNA__08275__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07588_ top.DUT.register\[19\]\[3\] net731 net727 top.DUT.register\[10\]\[3\] _02714_
+ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a221o_1
XANTENNA__10377__Y _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06539_ _01591_ _01631_ _01637_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__and3_4
X_09327_ top.pc\[16\] _04362_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or2_1
XANTENNA__09273__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07284__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09258_ net138 _04295_ _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08209_ _03173_ _03182_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__nand2_1
XANTENNA__09025__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ _04244_ _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__nor2_1
XANTENNA__09025__B2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_177_Right_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ net882 net884 top.a1.row2\[12\] _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and4b_1
XANTENNA__08304__A _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11151_ wb.curr_state\[0\] net855 _01434_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__o21a_1
XANTENNA__10045__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net1421 net251 net461 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
X_11082_ net917 net1300 net852 _05027_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__a31o_1
XANTENNA__08536__A0 _03456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ net259 net1884 net421 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__mux2_1
XANTENNA__09135__A _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13653__Q net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__B net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08839__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ _05843_ _05853_ _05841_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08839__B2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13723_ clknet_leaf_73_clk _01266_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10935_ top.a1.state\[2\] net893 vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ clknet_leaf_87_clk _01213_ net1008 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10866_ net1431 net155 net351 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12605_ clknet_leaf_104_clk _00169_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13585_ clknet_leaf_98_clk _01144_ net982 vssd1 vssd1 vccd1 vccd1 top.ramload\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10797_ net1451 net166 net447 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ clknet_leaf_93_clk _00100_ net999 vssd1 vssd1 vccd1 vccd1 top.pc\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07814__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ clknet_leaf_100_clk top.ru.next_FetchedInstr\[19\] net986 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07027__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _05229_ _05278_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__xnor2_1
X_12398_ clknet_leaf_89_clk _00034_ net1006 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ top.a1.dataIn\[25\] _05203_ _05211_ _05214_ _05218_ vssd1 vssd1 vccd1 vccd1
+ _05219_ sky130_fd_sc_hd__o41a_1
XFILLER_0_207_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11575__A top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_107_clk_X clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ clknet_leaf_52_clk _00583_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ top.DUT.register\[19\]\[22\] net633 net787 top.DUT.register\[3\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a22o_1
XANTENNA__10885__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06553__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08560_ net270 _03466_ _03472_ net274 vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07511_ top.a1.instruction\[16\] net524 _02637_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a21o_2
XFILLER_0_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08491_ net319 _03607_ _03597_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__o21ba_1
X_07442_ top.DUT.register\[19\]\[6\] net633 net787 top.DUT.register\[3\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07373_ top.DUT.register\[29\]\[7\] net701 net673 top.DUT.register\[16\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06324_ _01447_ _01461_ _01464_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__o21ai_1
X_09112_ _04168_ _04165_ _04028_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux2_1
XANTENNA__07266__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__X _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09043_ _04074_ _04097_ _04104_ _03728_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__or4b_1
X_06255_ net2354 top.ru.next_iready vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout309_A _02759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07018__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold410 top.DUT.register\[12\]\[22\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06186_ top.a1.halfData\[5\] _01414_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10373__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 top.DUT.register\[11\]\[31\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 top.DUT.register\[22\]\[19\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 top.DUT.register\[15\]\[15\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold454 top.DUT.register\[10\]\[22\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 top.DUT.register\[13\]\[25\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold476 top.DUT.register\[7\]\[6\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 top.DUT.register\[23\]\[4\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_2
Xhold498 top.DUT.register\[19\]\[16\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout912 _01408_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_2
X_09945_ net217 net1960 net433 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__mux2_1
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout580_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Left_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout934 net980 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_2
Xfanout945 net946 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_2
XANTENNA_fanout678_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07682__B _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__inv_2
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_2
Xhold1110 top.DUT.register\[5\]\[4\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
Xfanout989 net996 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_4
Xhold1121 top.DUT.register\[6\]\[17\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 top.pad.keyCode\[5\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08827_ _03192_ _03195_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nand2_1
Xhold1143 top.DUT.register\[10\]\[0\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 top.DUT.register\[20\]\[14\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06298__B net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 top.DUT.register\[26\]\[29\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 top.DUT.register\[22\]\[17\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 top.a1.row2\[15\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _02037_ _03091_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_142_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ top.DUT.register\[19\]\[1\] net634 net788 top.DUT.register\[3\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__a22o_1
X_08689_ _02951_ _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ net200 net2123 net383 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
XANTENNA__12910__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Left_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ net1902 net235 net450 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07257__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ net255 net1844 net386 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
X_13370_ clknet_leaf_18_clk _00934_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12321_ top.pad.count\[0\] net912 vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12252_ _01382_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__nand2_1
XANTENNA__08034__A _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12552__Q top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net1208 _05079_ _05088_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__a21o_1
X_12183_ _06050_ _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Left_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ net917 net1453 net852 _05053_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a31o_1
XANTENNA__08509__A0 _03426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A1 _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06783__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ net80 net864 net828 net1256 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a22o_1
XANTENNA__10503__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net205 net2155 net426 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_174_Left_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09485__A1 _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ _05797_ _05829_ _05830_ _05794_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12590__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13706_ clknet_leaf_75_clk _01254_ net1090 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06299__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ net180 net1856 net442 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ _05747_ _05749_ _05730_ _05733_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_67_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13637_ clknet_leaf_61_clk net1282 net1100 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09237__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10849_ net2179 net208 net351 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07248__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ clknet_leaf_84_clk _01127_ net1017 vssd1 vssd1 vccd1 vccd1 top.a1.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12519_ clknet_leaf_80_clk _00083_ net1002 vssd1 vssd1 vccd1 vccd1 top.pc\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13499_ clknet_leaf_48_clk _01063_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_183_Left_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08748__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13884__1134 vssd1 vssd1 vccd1 vccd1 _13884__1134/HI net1134 sky130_fd_sc_hd__conb_1
XANTENNA__07420__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06223__B2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 net210 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
Xfanout219 _04732_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10480__Y _04959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ top.DUT.register\[25\]\[31\] net773 net676 top.DUT.register\[18\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06774__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ top.pc\[13\] _04329_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__and2_1
X_06942_ top.DUT.register\[20\]\[21\] net579 net551 top.DUT.register\[24\]\[21\] _02068_
+ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__a221o_1
XANTENNA__10413__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ net794 _04682_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__or2_1
XANTENNA__09712__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ top.DUT.register\[22\]\[22\] net753 net688 top.DUT.register\[1\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ net280 _03679_ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__o21ai_1
X_09592_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08543_ net320 _03657_ _03655_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_173_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout161_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout259_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07487__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08474_ _02450_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08119__A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07425_ top.DUT.register\[10\]\[6\] net729 net677 top.DUT.register\[18\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1070_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout426_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07239__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ top.DUT.register\[2\]\[8\] net659 net611 top.DUT.register\[14\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06307_ net2199 _01445_ _01446_ net881 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07287_ top.DUT.register\[27\]\[9\] net776 net760 top.DUT.register\[26\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ net275 _03483_ _03741_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__o211a_1
X_06238_ net1707 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[14\] sky130_fd_sc_hd__and2_1
XANTENNA__06462__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold240 top.DUT.register\[28\]\[10\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_06169_ top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XANTENNA__08203__A2 _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 top.DUT.register\[28\]\[2\] vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 top.DUT.register\[27\]\[31\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 top.DUT.register\[14\]\[25\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07411__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 top.DUT.register\[28\]\[12\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 top.a1.data\[4\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout962_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _01527_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06765__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 _01522_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
XANTENNA__10323__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09928_ net150 net2286 net433 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__mux2_1
Xfanout742 _01519_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_4
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_8
Xfanout764 _01509_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout775 _01502_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
XANTENNA__09703__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout786 _01657_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_2
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _04853_ _04854_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__o21ai_2
Xfanout797 _04969_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08795__Y _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ clknet_leaf_25_clk _00434_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07190__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _05672_ _05676_ _05651_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07478__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__A1 top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ _05589_ _05600_ _05594_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09132__B _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08029__A _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10703_ net158 top.DUT.register\[24\]\[28\] net380 vssd1 vssd1 vccd1 vccd1 _00886_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11683_ _05494_ _05516_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_81_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13422_ clknet_leaf_118_clk _00986_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10634_ net175 net2289 net389 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13353_ clknet_leaf_2_clk _00917_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10565_ net211 net1734 net359 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ top.lcd.cnt_500hz\[9\] _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__or2_1
XANTENNA__07650__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13284_ clknet_leaf_42_clk _00848_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10496_ net182 net1278 net365 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12235_ top.lcd.cnt_20ms\[13\] top.lcd.cnt_20ms\[12\] top.lcd.cnt_20ms\[11\] top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or4bb_1
XANTENNA__07402__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _06026_ _06028_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06756__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ net49 net858 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__and2_1
X_12097_ _05953_ _05962_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_207_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08211__B net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ net2321 net855 _01432_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__o21a_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
XANTENNA__07705__A1 top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07181__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09458__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12999_ clknet_leaf_8_clk _00563_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07469__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11265__B2 top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07210_ top.DUT.register\[25\]\[15\] net772 net719 top.DUT.register\[2\]\[15\] _02336_
+ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08190_ net294 _02875_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__nand2_1
XANTENNA__12214__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08969__B1 _02947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ top.DUT.register\[31\]\[12\] net784 net628 top.DUT.register\[9\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_191_Left_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10408__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07641__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ top.a1.instruction\[4\] _01581_ _01488_ _01480_ vssd1 vssd1 vccd1 vccd1 _02199_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10143__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__B _02427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ _01860_ _03100_ _01821_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__a21o_1
XANTENNA__09932__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ net233 net1468 net438 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
X_06925_ top.DUT.register\[26\]\[21\] net762 net707 top.DUT.register\[15\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a22o_1
XANTENNA__09697__A1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout376_A _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ top.a1.halfData\[3\] _01472_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__or2_1
XANTENNA__07960__B _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06856_ top.DUT.register\[4\]\[23\] net767 net674 top.DUT.register\[18\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XANTENNA__07172__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09233__A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13751__Q top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ _04589_ _04592_ _04593_ _04607_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout543_A _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06787_ top.DUT.register\[27\]\[24\] net776 _01535_ top.DUT.register\[3\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ _02903_ _03574_ _02236_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09520__X _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ _02450_ _03573_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__xor2_2
XFILLER_0_148_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13261__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__A1 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ _02527_ _02529_ _02531_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__or4_1
XANTENNA__07880__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12205__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ _02588_ _03177_ net483 _02587_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07339_ top.DUT.register\[26\]\[8\] net759 net720 top.DUT.register\[14\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10350_ net1414 net200 net394 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06986__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _03752_ _03768_ _03790_ _03806_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ net2005 net207 net401 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _05884_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__or2_1
XANTENNA__10053__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09127__B _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 _01661_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_8
Xfanout561 _01650_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_4
Xfanout572 _01635_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_8
Xfanout583 _01513_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_4
Xfanout594 _04041_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_4
X_12922_ clknet_leaf_15_clk _00486_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07699__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08458__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08360__B2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ clknet_leaf_6_clk _00417_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13661__Q net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11804_ _05614_ _05635_ _05665_ _05613_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12784_ clknet_leaf_121_clk _00348_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13883__1133 vssd1 vssd1 vccd1 vccd1 _13883__1133/HI net1133 sky130_fd_sc_hd__conb_1
XFILLER_0_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11735_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08663__A2 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13373__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ _05507_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__nand2_2
X_13405_ clknet_leaf_112_clk _00969_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net244 top.DUT.register\[22\]\[6\] net391 vssd1 vssd1 vccd1 vccd1 _00800_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10228__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11597_ _05465_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07623__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ clknet_leaf_13_clk _00900_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10548_ net263 net1499 net358 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__06977__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ clknet_leaf_4_clk _00831_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10479_ net140 net1768 net371 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12218_ net1171 _06057_ net589 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
X_13198_ clknet_leaf_115_clk _00762_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06729__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ top.a1.dataIn\[2\] _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__xor2_2
XFILLER_0_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10898__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A1 _03437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__Y _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__B _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ top.DUT.register\[19\]\[26\] net733 net729 top.DUT.register\[10\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
X_07690_ top.DUT.register\[13\]\[0\] net678 _02812_ _02816_ vssd1 vssd1 vccd1 vccd1
+ _02817_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07154__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ _01760_ _01762_ _01764_ _01767_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06901__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _04404_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_121_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06572_ top.DUT.register\[28\]\[29\] net586 net698 top.DUT.register\[23\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ net468 _03415_ _03421_ net476 _03428_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ top.pc\[14\] _04325_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__and2_1
X_08242_ _03365_ _03366_ net302 vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07301__A _02427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ net292 _03054_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__nand2_1
XANTENNA__10138__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09480__A_N net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ top.DUT.register\[21\]\[12\] net693 _02237_ _02250_ vssd1 vssd1 vccd1 vccd1
+ _02251_ sky130_fd_sc_hd__a211o_1
XANTENNA__08968__A1_N _02989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06968__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07055_ top.DUT.register\[14\]\[10\] net721 net675 top.DUT.register\[18\]\[10\] _02181_
+ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1033_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13746__Q top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07971__A _01909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _03079_ _03082_ _02993_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout660_A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _01515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ net513 _02034_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__nor2_1
XANTENNA__10601__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ top.DUT.register\[19\]\[17\] net631 net785 top.DUT.register\[3\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__a22o_1
XANTENNA__07145__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09627_ _04650_ _04652_ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__or3b_1
X_06839_ top.DUT.register\[3\]\[23\] net785 _01965_ vssd1 vssd1 vccd1 vccd1 _01966_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09558_ _04579_ _04590_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08509_ _03426_ _03624_ net310 vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ _04501_ _04503_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__nand2_1
XANTENNA__08645__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11520_ _05321_ _05339_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07853__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _05311_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10048__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ net191 net2239 net330 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11382_ _05219_ _05225_ _05217_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06959__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ clknet_leaf_26_clk _00685_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ net2173 net146 net397 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_185_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07865__B _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__Y _03437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13157__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13052_ clknet_leaf_56_clk _00616_ net1086 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10264_ net1492 net147 net455 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__mux2_1
X_12003_ _05871_ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nand2_1
X_10195_ net156 top.DUT.register\[9\]\[28\] net411 vssd1 vssd1 vccd1 vccd1 _00406_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07384__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout380 _04949_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_13__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__06592__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout391 _04944_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11468__A1 top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06497__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07136__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12905_ clknet_leaf_3_clk _00469_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13885_ net1135 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12836_ clknet_leaf_40_clk _00400_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ clknet_leaf_114_clk _00331_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09833__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06647__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11718_ _05549_ _05571_ _05572_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12698_ clknet_leaf_16_clk _00262_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09046__C1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11649_ _05493_ _05499_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__xnor2_2
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12196__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold806 top.DUT.register\[4\]\[28\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold817 top.DUT.register\[15\]\[24\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold828 top.DUT.register\[15\]\[5\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_8_clk _00883_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold839 top.DUT.register\[17\]\[25\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12470__Q top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08860_ _03922_ _03958_ _01818_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_209_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07375__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ top.DUT.register\[28\]\[19\] net653 net605 top.DUT.register\[18\]\[19\] _02937_
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__a221o_1
X_08791_ net316 _03259_ _03559_ _03891_ net481 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o32a_2
XANTENNA__06583__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__C1 _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10421__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07742_ top.DUT.register\[1\]\[1\] net687 _02862_ _02868_ vssd1 vssd1 vccd1 vccd1
+ _02869_ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ top.DUT.register\[2\]\[0\] net659 net556 top.DUT.register\[6\]\[0\] _02799_
+ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08875__A2 _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ _04453_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__nand2b_1
X_06624_ top.DUT.register\[20\]\[28\] net749 net682 top.DUT.register\[7\]\[28\] _01750_
+ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09343_ _04388_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06555_ net900 _01592_ net801 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__and3b_4
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout241_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout339_A _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09230__B _02427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ net894 top.pc\[13\] _04293_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__and3_1
X_06486_ _01605_ _01612_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__or2_2
XFILLER_0_191_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08225_ net313 _03350_ _03328_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12187__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ _01755_ net297 vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08414__X _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07063__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _02184_ _02232_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08087_ _03212_ _03213_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07038_ _02163_ _02164_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_209_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13882__1132 vssd1 vssd1 vccd1 vccd1 _13882__1132/HI net1132 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_149_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _03332_ _03380_ _03452_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__and4_1
XANTENNA__06574__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__B2 _03438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ net844 _04977_ top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ clknet_leaf_84_clk _01229_ net1015 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10882_ net1611 net209 net347 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12621_ clknet_leaf_32_clk _00185_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__A2 _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07212__Y _02339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ clknet_leaf_69_clk _00116_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ _05349_ _05371_ _05338_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12483_ clknet_leaf_94_clk net34 net997 vssd1 vssd1 vccd1 vccd1 top.testpc.en_latched
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_191_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11434_ _05265_ _05291_ _05270_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_78_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06780__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11365_ _05233_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_100_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10506__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13104_ clknet_leaf_122_clk _00668_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10316_ net1969 net201 net399 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11296_ top.a1.row1\[109\] _05161_ _05166_ _05169_ _05170_ vssd1 vssd1 vccd1 vccd1
+ _05171_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08003__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13035_ clknet_leaf_30_clk _00599_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ net1397 net200 net456 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__mux2_1
XANTENNA__07357__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ net221 net1718 net411 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10241__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10113__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13868_ net1155 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_12819_ clknet_leaf_5_clk _00383_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13799_ clknet_leaf_65_clk _01342_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06340_ _01472_ vssd1 vssd1 vccd1 vccd1 top.edg2.button_i sky130_fd_sc_hd__inv_2
XANTENNA__09050__B _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12465__Q top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06271_ top.ramload\[15\] net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[15\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_72_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08010_ top.DUT.register\[3\]\[31\] net788 net784 top.DUT.register\[31\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a22o_1
Xhold603 top.DUT.register\[21\]\[2\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 top.DUT.register\[11\]\[7\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10416__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold625 top.DUT.register\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 top.DUT.register\[31\]\[14\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 top.DUT.register\[10\]\[26\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold658 top.DUT.register\[30\]\[20\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _04676_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__nor2_2
XFILLER_0_122_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold669 top.ramload\[8\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08888__Y _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ net519 _04006_ _04008_ _04005_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__o211a_1
X_09892_ _04578_ net527 net333 top.a1.dataIn\[28\] net335 vssd1 vssd1 vccd1 vccd1
+ _04887_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07348__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09506__A _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _01821_ _01860_ _03100_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__nand3_1
XANTENNA__10352__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06556__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10151__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ _03545_ _03745_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__nand2_2
XANTENNA__09940__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07725_ top.DUT.register\[30\]\[1\] net617 net542 top.DUT.register\[22\]\[1\] _02851_
+ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_69_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout456_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _02781_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__nand2_2
XFILLER_0_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07520__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ _01713_ _01732_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout623_A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ top.DUT.register\[11\]\[3\] net755 net735 top.DUT.register\[24\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08128__Y _03255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09326_ top.pc\[16\] _04362_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06538_ _01628_ _01631_ _01634_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__and3_4
XANTENNA__07808__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ net134 _04301_ _04308_ _04309_ net911 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06469_ top.a1.instruction\[13\] net901 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08208_ _03156_ _03160_ _03173_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__and3_4
X_09188_ top.pc\[7\] _02567_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ _01929_ net292 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10326__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07587__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ net897 net1602 _05059_ _05062_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ net1506 net257 net462 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ net40 net861 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07339__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ net265 net1490 net423 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__mux2_1
XANTENNA__06547__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10061__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _05825_ _05845_ _05840_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13722_ clknet_leaf_73_clk _01265_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10934_ net140 net1915 net444 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09151__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13653_ clknet_leaf_86_clk _01212_ net1014 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10865_ net2068 net157 net352 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12604_ clknet_leaf_55_clk _00168_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13584_ clknet_leaf_97_clk _01143_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10796_ net1500 net170 net446 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12535_ clknet_leaf_90_clk _00099_ net998 vssd1 vssd1 vccd1 vccd1 top.pc\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[18\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[18\] sky130_fd_sc_hd__dfrtp_4
X_11417_ _05285_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ clknet_leaf_88_clk _00033_ net1005 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08775__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ top.a1.dataIn\[27\] _05196_ _05198_ _05201_ vssd1 vssd1 vccd1 vccd1 _05218_
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11279_ _05098_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__nor2_1
XANTENNA__09724__B1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ clknet_leaf_51_clk _00582_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ top.a1.instruction\[11\] _01477_ _01620_ net900 vssd1 vssd1 vccd1 vccd1 _02637_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ net312 _03372_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09061__A _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07441_ top.DUT.register\[17\]\[6\] net646 net610 top.DUT.register\[12\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06710__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881__1131 vssd1 vssd1 vccd1 vccd1 _13881__1131/HI net1131 sky130_fd_sc_hd__conb_1
X_07372_ top.DUT.register\[22\]\[7\] net751 net667 top.DUT.register\[5\]\[7\] _02498_
+ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09111_ _04170_ _04154_ _04145_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__mux2_1
X_06323_ _01333_ _01459_ _01463_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__or3_1
XFILLER_0_174_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11062__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09042_ _03598_ _03828_ _04098_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06254_ net1362 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[30\] sky130_fd_sc_hd__and2_1
XFILLER_0_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 top.DUT.register\[12\]\[5\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10146__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06185_ top.a1.halfData\[1\] top.a1.halfData\[2\] top.a1.halfData\[3\] vssd1 vssd1
+ vccd1 vccd1 _01414_ sky130_fd_sc_hd__nand3b_1
Xhold411 top.DUT.register\[9\]\[9\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 top.DUT.register\[12\]\[1\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07569__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 top.DUT.register\[5\]\[31\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 top.DUT.register\[15\]\[11\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 top.DUT.register\[20\]\[21\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 top.DUT.register\[29\]\[27\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 top.DUT.register\[20\]\[3\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout902 top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_2
X_09944_ net227 net2197 net434 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__mux2_1
Xhold488 top.DUT.register\[30\]\[25\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 top.DUT.register\[22\]\[1\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout924 net934 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_55_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09715__B1 _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net980 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08140__A _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06212__X _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ top.pc\[27\] _04557_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
Xfanout957 net964 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_2
XANTENNA__13754__Q top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout968 net979 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_2
Xhold1100 top.DUT.register\[5\]\[24\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout573_A _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1111 top.DUT.register\[9\]\[17\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net980 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ net305 _03857_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__or2_1
Xhold1122 top.DUT.register\[18\]\[28\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 top.DUT.register\[30\]\[18\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 top.DUT.register\[15\]\[23\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 top.DUT.register\[22\]\[12\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 top.DUT.register\[11\]\[6\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1177 top.DUT.register\[27\]\[20\] vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net478 _03852_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21boi_4
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 top.DUT.register\[28\]\[31\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07708_ _01616_ _02833_ _02834_ _02832_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__a31o_2
X_08688_ _02993_ _03779_ _02991_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07639_ top.DUT.register\[14\]\[2\] net720 net716 top.DUT.register\[2\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06701__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12539__RESET_B net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ net1976 net241 net450 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09309_ _04344_ _04345_ _04346_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_192_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10581_ net261 net1763 net385 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XANTENNA__08454__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12320_ top.pad.count\[0\] net912 vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ net1187 _06064_ _06078_ net1108 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__o211a_1
XANTENNA__10056__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08034__B _03155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08757__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ net851 _05074_ _05078_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__and3_1
X_12182_ _06039_ _06044_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__a21boi_2
XANTENNA__06768__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11133_ net58 net857 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__and2_1
XANTENNA__07365__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11108__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__B1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net79 net858 net829 net1177 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__a22o_1
XANTENNA__09182__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net213 net2328 net427 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XANTENNA__08985__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07732__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06940__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11966_ _05831_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06299__A2 _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ net195 net1796 net444 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
X_13705_ clknet_leaf_75_clk _01253_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11897_ _05717_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13636_ clknet_leaf_61_clk net1199 net1102 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10848_ net1735 net219 net351 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13567_ clknet_leaf_84_clk _01126_ net1017 vssd1 vssd1 vccd1 vccd1 top.a1.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ net1504 net238 net445 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ clknet_leaf_70_clk top.a1.nextHex\[7\] net1103 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13498_ clknet_leaf_18_clk _01062_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12449_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[1\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06759__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13750__RESET_B net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlymetal6s2s_1
X_07990_ _03113_ _03115_ _03116_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06941_ top.DUT.register\[13\]\[21\] net650 net646 top.DUT.register\[17\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a22o_1
X_09660_ net794 _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__nor2_1
X_06872_ top.DUT.register\[25\]\[22\] net773 net722 top.DUT.register\[14\]\[22\] _01998_
+ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a221o_1
XANTENNA__07184__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ net288 _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__or2_1
XANTENNA__07723__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ net910 _04169_ _04180_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and3_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06931__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _03409_ _03545_ _03654_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nand3_1
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _02493_ _03555_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07424_ top.DUT.register\[27\]\[6\] net778 net587 top.DUT.register\[28\]\[6\] _02550_
+ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07355_ top.DUT.register\[19\]\[8\] net631 net781 top.DUT.register\[31\]\[8\] _02481_
+ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout321_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout419_A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06306_ top.lcd.currentState\[0\] net885 net824 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07286_ _02408_ _02410_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__or3_1
XANTENNA__06998__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13749__Q top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09025_ net275 _03495_ _03719_ net313 _03256_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06237_ net1320 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[13\] sky130_fd_sc_hd__and2_1
XFILLER_0_131_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold230 top.DUT.register\[11\]\[16\] vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 top.a1.hexop\[2\] vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold252 top.DUT.register\[29\]\[5\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 top.DUT.register\[13\]\[24\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 top.DUT.register\[17\]\[14\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 top.DUT.register\[14\]\[29\] vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 top.DUT.register\[11\]\[17\] vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_4
Xfanout721 _01527_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
Xfanout732 _01522_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
X_09927_ net464 _04917_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nand2_4
Xfanout743 _01518_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 _01516_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_4
Xfanout765 _01509_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 _01502_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_4
X_09858_ net833 _04517_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__o21ba_1
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_4
XANTENNA__07175__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout798 _04969_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_198_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07714__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__B2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ net268 _03742_ _03771_ _03578_ _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ net802 _04790_ _04791_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a31o_1
XANTENNA__06922__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11820_ _05641_ _05646_ _05672_ _05676_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_1_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _05603_ _05620_ _05617_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08029__B _03155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ net161 net1958 net378 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
X_11682_ _05532_ _05539_ _05546_ _05548_ _05550_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13421_ clknet_leaf_32_clk _00985_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ net183 net1919 net392 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_34_clk _00916_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10564_ net215 net2322 net357 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08045__A _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13659__Q net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _06109_ net588 _06108_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__and3b_1
X_13283_ clknet_leaf_50_clk _00847_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10495_ net197 net2084 net367 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__mux2_1
X_12234_ top.lcd.cnt_20ms\[9\] top.lcd.cnt_20ms\[7\] top.lcd.cnt_20ms\[6\] top.lcd.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__or4b_1
XFILLER_0_20_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13533__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10514__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _06030_ _06033_ _06027_ _06029_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net918 net1328 net855 _05044_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a31o_1
X_12096_ _05965_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_207_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ net1182 net856 net825 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__a21o_1
XANTENNA__07166__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06913__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12998_ clknet_leaf_9_clk _00562_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11291__D net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _05754_ _05786_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_139_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13619_ clknet_leaf_45_clk net1207 net1081 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07778__B _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08969__B2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ top.DUT.register\[19\]\[12\] net634 net788 top.DUT.register\[3\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12473__Q top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07071_ _02193_ _02197_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10424__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07944__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ _01865_ _03099_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__or2_1
X_09712_ _03593_ net340 net336 _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__o211a_1
X_06924_ top.DUT.register\[27\]\[21\] net777 net757 top.DUT.register\[11\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a22o_1
XANTENNA__07157__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09697__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _04646_ _04647_ _01472_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__o21ai_1
X_06855_ _01976_ _01978_ _01980_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06904__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout369_A _04958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09574_ _04589_ _04592_ _04593_ _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__or4_1
XANTENNA__09233__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06786_ _01911_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10379__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08525_ net1306 net837 net816 _03640_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout536_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08456_ _02450_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08417__X _03537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07407_ top.DUT.register\[20\]\[7\] net576 net630 top.DUT.register\[9\]\[7\] _02533_
+ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a221o_1
XANTENNA__12205__A1 top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ net269 _03507_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nand2_1
XANTENNA__06683__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__B2 top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10216__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ top.DUT.register\[17\]\[8\] net726 net692 top.DUT.register\[21\]\[8\] _02464_
+ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07632__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ top.DUT.register\[25\]\[14\] net625 net617 top.DUT.register\[30\]\[14\] _02384_
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a221o_1
X_09008_ _03827_ _03843_ _03860_ _03875_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__nand4b_1
X_10280_ net2214 net221 net403 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10334__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__A1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _01671_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout551 _01661_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_4
XANTENNA__09137__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_8
Xfanout573 _01635_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_4
Xfanout584 _01512_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 _01670_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_8
X_12921_ clknet_leaf_37_clk _00485_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06400__X _01527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12852_ clknet_leaf_45_clk _00416_ net1080 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11803_ _05660_ _05668_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_14_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08648__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12783_ clknet_leaf_20_clk _00347_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08982__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11734_ _05589_ _05599_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__nor2_2
XFILLER_0_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07320__A0 _02427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11665_ _05517_ _05518_ _05521_ _05504_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__o31a_1
XANTENNA__06674__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10509__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ net248 net1817 net390 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__mux2_1
X_13404_ clknet_leaf_54_clk _00968_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ _05430_ _05453_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13335_ clknet_leaf_105_clk _00899_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10547_ net148 top.DUT.register\[20\]\[0\] net357 vssd1 vssd1 vccd1 vccd1 _00730_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07885__Y _03012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ clknet_leaf_48_clk _00830_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_23_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10478_ net146 net1812 net370 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12217_ net1170 _06056_ net590 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XANTENNA__10244__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ clknet_leaf_32_clk _00761_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07387__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _06013_ _06017_ _06011_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ _05947_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__nand2_1
XANTENNA__07139__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06640_ top.DUT.register\[20\]\[28\] net578 _01758_ _01765_ _01766_ vssd1 vssd1 vccd1
+ vccd1 _01767_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_189_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06571_ top.DUT.register\[2\]\[29\] net717 net676 top.DUT.register\[18\]\[29\] _01696_
+ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08310_ net483 _03413_ _03433_ net479 _03427_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09290_ net911 top.pc\[13\] _04340_ net899 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__o211a_1
XANTENNA__06693__A _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _03210_ _03214_ net276 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06665__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10419__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12199__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08172_ _02339_ net297 vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ top.DUT.register\[1\]\[12\] net686 net684 top.DUT.register\[7\]\[12\] _02249_
+ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_41_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13083__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__S net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ top.DUT.register\[4\]\[10\] net770 net760 top.DUT.register\[26\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a22o_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__07090__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA__13012__RESET_B net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08492__A1_N _03183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__B _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A _03179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _03079_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nand2_1
X_06907_ net808 _02033_ _01625_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__o21a_1
X_07887_ top.DUT.register\[8\]\[17\] net568 net540 top.DUT.register\[22\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_50_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08878__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ _04646_ _04647_ _04648_ _04645_ _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__o221a_1
X_06838_ top.DUT.register\[31\]\[23\] net781 net779 top.DUT.register\[15\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
XANTENNA__07550__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ _04575_ _04581_ _04590_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__B _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06769_ top.DUT.register\[15\]\[25\] _01655_ net782 top.DUT.register\[31\]\[25\]
+ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_35_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ _03536_ _03623_ net307 vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09488_ _04525_ _04526_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07302__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ _03219_ net272 _03253_ net268 vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a22o_1
XANTENNA__10329__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06656__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ _05309_ _05280_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__and2b_1
XFILLER_0_163_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10401_ net203 net2000 net330 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
X_11381_ _05249_ _05250_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13120_ clknet_leaf_43_clk _00684_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ net1697 net152 net398 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__mux2_1
XANTENNA__09419__A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_185_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13051_ clknet_leaf_58_clk _00615_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10263_ net1495 net153 net456 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08042__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12002_ _05843_ _05853_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__xor2_1
X_10194_ net163 net1939 net409 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 _04958_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_4
Xfanout381 _04947_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_6
Xfanout392 _04944_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_4
XFILLER_0_205_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12904_ clknet_leaf_35_clk _00468_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13884_ net1134 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_186_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07541__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06895__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12835_ clknet_leaf_33_clk _00399_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__C1 _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ clknet_leaf_14_clk _00330_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10979__A1 top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11717_ _05549_ _05572_ _05571_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06647__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ clknet_leaf_36_clk _00261_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10239__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09046__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11648_ _05500_ _05515_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11859__A top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_2
X_11579_ _05439_ _05448_ _05441_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold807 top.DUT.register\[22\]\[28\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold818 top.DUT.register\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_9_clk _00882_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 top.DUT.register\[27\]\[0\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13101__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_208_Right_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ clknet_leaf_26_clk _00813_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07810_ top.DUT.register\[17\]\[19\] net645 net602 top.DUT.register\[10\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a22o_1
XANTENNA__08572__A2 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13251__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ _01953_ net470 _03878_ net478 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a22o_1
X_07741_ top.DUT.register\[24\]\[1\] net737 net734 top.DUT.register\[19\]\[1\] _02861_
+ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07672_ top.DUT.register\[1\]\[0\] net655 net548 top.DUT.register\[24\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__a22o_1
XANTENNA__07532__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ top.pc\[21\] _04443_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__nand2_1
X_06623_ top.DUT.register\[30\]\[28\] net715 _01737_ _01746_ vssd1 vssd1 vccd1 vccd1
+ _01750_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06694__Y _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ top.pc\[17\] _04379_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06554_ top.DUT.register\[21\]\[30\] net572 net648 top.DUT.register\[13\]\[30\] _01680_
+ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08408__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06638__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ net911 net894 _04324_ net899 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06485_ _01578_ _01582_ _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10149__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08224_ net283 _03349_ _03281_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__a21o_2
XANTENNA__09938__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__Y _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08155_ net285 _03279_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout401_A _04939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07599__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ _02184_ _02232_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__or2_1
XANTENNA__08260__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ net289 _02928_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08143__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07037_ _02142_ _02162_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06810__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__S net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ _03171_ net476 vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nor2_1
X_07939_ top.DUT.register\[15\]\[16\] net780 _03055_ _03065_ vssd1 vssd1 vccd1 vccd1
+ _03066_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ net2126 _04980_ _04979_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_162_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09609_ _04628_ net851 _04637_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a21o_1
XANTENNA__06877__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ net1664 net220 net348 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12620_ clknet_leaf_10_clk _00184_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09758__A1_N _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06629__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ clknet_leaf_71_clk _00115_ net1093 vssd1 vssd1 vccd1 vccd1 top.a1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10059__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _05349_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12482_ clknet_leaf_69_clk _00050_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.debounce
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11433_ _05289_ _05290_ _05264_ _05271_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_78_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11364_ top.a1.dataIn\[19\] _05223_ _05224_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__and3_1
XANTENNA__07054__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12987__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10315_ net1428 net209 net398 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
X_13103_ clknet_leaf_51_clk _00667_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ top.a1.row1\[13\] _05093_ _05097_ _05112_ top.a1.row1\[61\] vssd1 vssd1 vccd1
+ vccd1 _05170_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_210_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11138__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A _03171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ clknet_leaf_34_clk _00598_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10246_ net1544 net209 net456 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__mux2_1
Xfanout1110 net39 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_4
XANTENNA__08554__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ net226 net2140 net409 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09503__A1 top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13867_ net1154 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_159_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12818_ clknet_leaf_50_clk _00382_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ clknet_leaf_67_clk _01341_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12749_ clknet_leaf_23_clk _00313_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06270_ net1707 net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[14\] sky130_fd_sc_hd__and2_1
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07293__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold604 top.DUT.register\[16\]\[21\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 top.DUT.register\[26\]\[15\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold626 top.ramaddr\[15\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold637 top.DUT.register\[2\]\[25\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold648 top.DUT.register\[7\]\[26\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09960_ _01601_ _04678_ _04675_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__or3b_2
Xhold659 top.DUT.register\[30\]\[5\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08911_ _01693_ net487 _03694_ _03771_ _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__o221a_1
X_09891_ _04883_ _04884_ _01586_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08545__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10432__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ _01821_ _03941_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_191_Right_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08773_ _01992_ net487 net468 _01994_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__o221a_1
XANTENNA__06211__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07724_ top.DUT.register\[1\]\[1\] net657 net550 top.DUT.register\[24\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06308__B2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__A _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06859__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _02759_ net495 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout351_A _04963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06865__B _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _01713_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nand2b_1
X_07586_ top.DUT.register\[31\]\[3\] net743 net667 top.DUT.register\[5\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09325_ top.pc\[15\] _04349_ _04359_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__a21o_1
X_06537_ _01591_ net789 _01637_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__and3_4
XANTENNA__11065__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09256_ _04302_ _04307_ _01619_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_4_10__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ net902 net901 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__and2_1
XANTENNA__07284__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08207_ _02831_ _02880_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09187_ top.pc\[7\] _02567_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__nor2_1
XANTENNA__10607__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06399_ top.DUT.register\[31\]\[30\] net744 _01520_ top.DUT.register\[17\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08138_ net1300 net839 _03263_ net815 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08069_ _03194_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10100_ net2248 net259 net459 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__mux2_1
XANTENNA__07992__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ net97 net862 net826 net1233 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ net151 net1620 net421 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10342__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__D _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__Y _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11982_ _05849_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__and2_1
X_13721_ clknet_leaf_67_clk _00004_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10933_ net144 net1880 net442 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13652_ clknet_leaf_87_clk _01211_ net1008 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
X_10864_ net1626 net161 net349 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13115__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ clknet_leaf_59_clk _00167_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13583_ clknet_leaf_98_clk _01142_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10795_ net1701 net171 net446 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12534_ clknet_leaf_90_clk _00098_ net998 vssd1 vssd1 vccd1 vccd1 top.pc\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06483__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ clknet_leaf_97_clk top.ru.next_FetchedInstr\[17\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10517__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07027__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08224__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _05253_ _05284_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__or2_1
X_12396_ clknet_leaf_88_clk _00032_ net1006 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12664__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11347_ _05182_ _05197_ _05216_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07983__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _05105_ _05112_ _05153_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or4_1
XANTENNA__08511__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10229_ net158 net2253 net408 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__mux2_1
X_13017_ clknet_leaf_36_clk _00581_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09724__B2 top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10252__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1 top.ramstore\[12\] vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07440_ _02566_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12476__Q top.a1.instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07371_ top.DUT.register\[27\]\[7\] net776 net767 top.DUT.register\[4\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__a22o_1
XANTENNA__06972__Y _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09110_ _04169_ _04171_ net895 vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__a21oi_1
X_06322_ _01451_ _01452_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_118_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07266__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09041_ _03964_ _04067_ _04100_ _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_40_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06253_ net1363 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[29\] sky130_fd_sc_hd__and2_1
XFILLER_0_154_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10427__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07018__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06184_ top.a1.halfData\[3\] _01412_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold401 top.DUT.register\[1\]\[24\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold412 top.DUT.register\[21\]\[18\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 top.DUT.register\[12\]\[29\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10373__D net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold434 top.DUT.register\[1\]\[25\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 top.DUT.register\[19\]\[21\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold456 top.DUT.register\[7\]\[10\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 top.DUT.register\[16\]\[7\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__B1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 top.DUT.register\[5\]\[13\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 top.DUT.register\[31\]\[2\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ net181 net2043 net433 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__mux2_1
XANTENNA__08421__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout903 top.a1.instruction\[12\] vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
XFILLER_0_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net916 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
Xfanout925 net933 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10162__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout947 net955 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
X_09874_ top.pc\[27\] _04557_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_1
Xfanout958 net964 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_4
Xhold1101 top.a1.hexop\[3\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07037__A _02142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 top.DUT.register\[2\]\[5\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1123 top.DUT.register\[15\]\[10\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _03100_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__nand2_1
Xhold1134 top.DUT.register\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 top.DUT.register\[9\]\[3\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 top.DUT.register\[16\]\[0\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1167 top.a1.row2\[25\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _03511_ _03771_ _03860_ _03184_ _03854_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__o221a_1
Xhold1178 top.DUT.register\[13\]\[23\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 top.DUT.register\[21\]\[8\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09252__A _02142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07707_ _02206_ _02785_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ net1262 net838 net818 _03795_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ top.DUT.register\[1\]\[2\] net685 net681 top.DUT.register\[7\]\[2\] _02764_
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout900_A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ top.DUT.register\[23\]\[3\] net560 net603 top.DUT.register\[18\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09308_ top.pc\[15\] _04349_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07257__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10580_ net264 net2103 net388 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XANTENNA__08454__B2 _03572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10261__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10337__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09239_ net911 top.pc\[10\] _04292_ net899 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_9__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ _06065_ _06070_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ net1954 _05079_ _04636_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_170_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08034__C _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11210__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _06019_ _06031_ _06040_ _06042_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ net914 net1342 net855 _05052_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a31o_1
Xhold990 top.DUT.register\[2\]\[28\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10072__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__B2 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ net78 net864 net828 net1276 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__a22o_1
XANTENNA__07717__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net215 top.DUT.register\[4\]\[17\] net425 vssd1 vssd1 vccd1 vccd1 _00235_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09861__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__B _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10800__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11965_ _05752_ _05799_ _05832_ _05833_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__and4b_1
XANTENNA__13462__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_74_clk _01252_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ net199 net2114 net444 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
XANTENNA__07496__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net129 _05749_ _05764_ _05720_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a211o_1
X_13635_ clknet_leaf_114_clk net1218 net940 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net1589 net223 net349 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07248__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13566_ clknet_leaf_75_clk _01125_ net1088 vssd1 vssd1 vccd1 vccd1 top.a1.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ net1708 net240 net446 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__mux2_1
X_12517_ clknet_leaf_70_clk _00009_ net1103 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10247__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13497_ clknet_leaf_36_clk _01061_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[0\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12379_ _01483_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__inv_2
XANTENNA__07420__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06940_ top.DUT.register\[15\]\[21\] _01655_ net633 top.DUT.register\[19\]\[21\]
+ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06871_ top.DUT.register\[8\]\[22\] net742 net669 top.DUT.register\[5\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08610_ _03298_ _03302_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10710__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09590_ top.pc\[31\] _04602_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_50_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08541_ net314 _03654_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_141_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09330__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ _03588_ _03589_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__nor2_1
XANTENNA__08684__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07423_ top.DUT.register\[3\]\[6\] net691 net670 top.DUT.register\[5\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XANTENNA__06695__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout147_A _04908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07354_ top.DUT.register\[3\]\[8\] net785 net779 top.DUT.register\[15\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07239__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06305_ _01447_ _01334_ _01335_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07285_ top.DUT.register\[12\]\[9\] net581 net721 top.DUT.register\[14\]\[9\] _02411_
+ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a221o_1
XANTENNA__10157__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _03891_ _03907_ _03931_ _03949_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout1056_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09946__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06236_ net1287 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[12\] sky130_fd_sc_hd__and2_1
XFILLER_0_198_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08703__X _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 top.DUT.register\[3\]\[24\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
Xhold231 top.DUT.register\[23\]\[1\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08422__Y _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 top.DUT.register\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 top.DUT.register\[30\]\[1\] vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07411__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 top.DUT.register\[7\]\[16\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 top.DUT.register\[19\]\[4\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _01536_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold297 top.DUT.register\[19\]\[19\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _01532_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_8
Xfanout722 net723 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
X_09926_ _04678_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__nor2_2
Xfanout733 net734 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 _01518_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1109_X net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout755 _01515_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_4
Xfanout766 _01509_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
X_09857_ _04518_ net527 net332 top.a1.dataIn\[25\] net334 vssd1 vssd1 vccd1 vccd1
+ _04855_ sky130_fd_sc_hd__a221o_1
Xfanout777 _01502_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
Xfanout788 _01657_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XANTENNA_fanout948_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13460__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13485__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10620__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _01908_ net485 _03909_ _01907_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_198_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09788_ top.a1.dataIn\[18\] net332 _04792_ net334 vssd1 vssd1 vccd1 vccd1 _04793_
+ sky130_fd_sc_hd__a211o_1
X_08739_ _03837_ _03838_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09321__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ top.a1.dataIn\[8\] _05602_ _05618_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__or3_1
XANTENNA__07478__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06686__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ net166 net2224 net380 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ _05548_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__and2_1
XFILLER_0_193_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ clknet_leaf_8_clk _00984_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10632_ net187 net1905 net392 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__mux2_1
XANTENNA__08427__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12223__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__A _02685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10067__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13351_ clknet_leaf_6_clk _00915_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10563_ net230 net2133 net360 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08045__B _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12302_ top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[8\] _06106_ vssd1 vssd1 vccd1 vccd1
+ _06109_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ clknet_leaf_41_clk _00846_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07650__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10494_ net199 net1607 net367 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__mux2_1
X_12233_ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07938__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__inv_2
XANTENNA__08061__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13675__Q top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ net48 net861 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__and2_1
XANTENNA__06610__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ _05949_ _05963_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_207_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11046_ net918 _01401_ wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_207_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10530__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__B net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12997_ clknet_leaf_119_clk _00561_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11948_ _05784_ _05786_ _05763_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07469__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06677__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11879_ _05705_ _05711_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a21o_2
XFILLER_0_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08792__C_N _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ clknet_leaf_82_clk net1186 net1012 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12214__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06429__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13549_ clknet_leaf_23_clk _01113_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07070_ _01478_ _01481_ _01576_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__o31a_1
XFILLER_0_152_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13358__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07641__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10705__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07929__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06601__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ net517 _01906_ _03098_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09554__A_N _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ top.pc\[9\] net803 _04718_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a211o_1
X_06923_ _02047_ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__or2_1
X_09642_ _04644_ _04651_ _04643_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10440__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ top.DUT.register\[28\]\[23\] net584 net689 top.DUT.register\[3\]\[23\] _01974_
+ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ _01560_ _04605_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__xnor2_1
X_06785_ top.DUT.register\[17\]\[24\] _01520_ net736 top.DUT.register\[24\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XANTENNA__10379__C net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ net888 top.pc\[11\] net538 _03639_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a22o_1
XANTENNA__08657__B2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06668__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ _02496_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout431_A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07406_ top.DUT.register\[2\]\[7\] net659 net782 top.DUT.register\[31\]\[7\] _02532_
+ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a221o_1
X_08386_ _03385_ _03506_ net305 vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08146__A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07337_ top.DUT.register\[25\]\[8\] net771 net671 top.DUT.register\[16\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09676__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07093__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ _02386_ _02388_ _02390_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__or4_1
XANTENNA__07632__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _03656_ _03676_ _03695_ _03720_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__and4_1
X_06219_ wb.curr_state\[0\] _01433_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06840__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ top.DUT.register\[17\]\[15\] _01520_ net732 top.DUT.register\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_187_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__C1 _04794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 _05079_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_4
Xfanout541 _01671_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_2
Xfanout552 net555 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_8
X_09909_ top.pc\[30\] _04605_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__xnor2_1
Xfanout563 _01650_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_4
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_4
Xfanout585 _01512_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_2
XANTENNA__10350__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ clknet_leaf_109_clk _00484_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout596 _01670_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07699__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12851_ clknet_leaf_5_clk _00415_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11802_ _05653_ _05657_ _05670_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12782_ clknet_leaf_116_clk _00346_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06659__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ _05560_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11664_ _05503_ _05523_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__xor2_2
XANTENNA__07871__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ clknet_leaf_52_clk _00967_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10615_ net253 net2018 net391 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__mux2_1
X_11595_ _05419_ _05464_ _05463_ _05423_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a2bb2o_2
X_13334_ clknet_leaf_121_clk _00898_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07623__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ net466 _04922_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06831__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10525__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13265_ clknet_leaf_3_clk _00829_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10477_ net153 net1922 net371 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12216_ net1169 top.a1.dataIn\[0\] net590 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13196_ clknet_leaf_11_clk _00760_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _06007_ _06004_ _06005_ _06015_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12078_ _05929_ _05946_ _05926_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10260__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ net8 net841 net811 net2251 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__o22a_1
XANTENNA__08887__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06898__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06570_ top.DUT.register\[30\]\[29\] net714 net669 top.DUT.register\[5\]\[29\] _01695_
+ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _03196_ _03207_ net276 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ net284 _03295_ _03281_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07122_ top.DUT.register\[31\]\[12\] net744 net720 top.DUT.register\[14\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XANTENNA__08253__X _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ top.DUT.register\[19\]\[10\] net731 net712 top.DUT.register\[30\]\[10\] _02179_
+ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a221o_1
XANTENNA__06822__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__09367__A2 top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06214__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1019_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _03035_ _03081_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout381_A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08327__B1 _02685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A _03255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ _02029_ _02031_ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nor3_4
XANTENNA__10170__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ top.DUT.register\[1\]\[17\] net655 net599 top.DUT.register\[10\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a22o_1
XANTENNA__06889__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ _04643_ _04651_ _04653_ _04644_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__o22a_1
X_06837_ top.DUT.register\[13\]\[23\] net647 net623 top.DUT.register\[25\]\[23\] _01963_
+ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout646_A _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _04579_ _04582_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__nor3_1
XFILLER_0_194_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06768_ top.DUT.register\[19\]\[25\] net632 net786 top.DUT.register\[3\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08507_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__inv_2
X_06699_ top.DUT.register\[12\]\[26\] net582 net758 top.DUT.register\[11\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
X_09487_ top.pc\[25\] _04508_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08438_ _03555_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nand2_1
XANTENNA__07853__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ net887 top.pc\[5\] net536 _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10400_ net211 net2161 net329 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__mux2_1
X_11380_ _05220_ _05225_ _05221_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08604__A _02401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10331_ net2266 net156 net399 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__mux2_1
XANTENNA__06813__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ net1887 net159 net457 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ clknet_leaf_21_clk _00614_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12001_ _05807_ _05870_ _05866_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__mux2_1
X_10193_ net166 net2096 net411 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09435__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout360 _04961_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_6
XFILLER_0_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout371 _04958_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06592__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10080__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout382 _04947_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_4
Xfanout393 net396 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
X_12903_ clknet_leaf_27_clk _00467_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13883_ net1133 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_201_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08993__B _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12834_ clknet_leaf_50_clk _00398_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12765_ clknet_leaf_108_clk _00329_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08057__Y _03184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11716_ _05574_ _05576_ _05581_ _05585_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ clknet_leaf_107_clk _00260_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ _05500_ _05504_ _05508_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__and3b_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 gpio_in[15] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
X_11578_ _05436_ _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold808 top.DUT.register\[6\]\[26\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
X_13317_ clknet_leaf_117_clk _00881_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap516 net517 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_2
XANTENNA__10255__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10529_ net1516 net180 net362 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__mux2_1
Xhold819 top.DUT.register\[7\]\[19\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ clknet_leaf_44_clk _00812_ net1082 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11156__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13179_ clknet_leaf_56_clk _00743_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06583__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07740_ _02858_ _02860_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__or3_1
XANTENNA__12479__Q top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07671_ top.DUT.register\[30\]\[0\] net615 net599 top.DUT.register\[10\]\[0\] _02797_
+ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__a221o_1
X_09410_ top.pc\[21\] _04443_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06622_ _01739_ _01741_ _01745_ _01748_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__or4_2
XFILLER_0_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09341_ top.pc\[17\] _04379_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__nor2_1
X_06553_ top.DUT.register\[7\]\[30\] net555 net616 top.DUT.register\[30\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_188_Left_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06484_ top.a1.instruction\[13\] _01489_ _01581_ _01610_ vssd1 vssd1 vccd1 vccd1
+ _01611_ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09272_ net134 _04317_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07835__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08223_ _03288_ _03348_ net299 vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout227_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08154_ _03279_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08424__A _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08796__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ _02212_ _02231_ net807 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_2
X_08085_ net295 _02970_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06215__Y _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07036_ _02142_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__nor2_1
XANTENNA__09954__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__X _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout596_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A2 _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout763_A _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _04045_ _04048_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06574__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ top.DUT.register\[31\]\[16\] net782 net600 top.DUT.register\[10\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ top.DUT.register\[25\]\[17\] net771 net747 top.DUT.register\[20\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout930_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__inv_2
X_10880_ net2163 net223 net345 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08981__A2_N net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09539_ _04558_ _04562_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10200__Y _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07287__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ clknet_leaf_71_clk _00114_ net1095 vssd1 vssd1 vccd1 vccd1 top.a1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07826__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _05364_ _05369_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a21o_2
X_12481_ clknet_leaf_95_clk top.ru.next_read_i net987 vssd1 vssd1 vccd1 vccd1 top.Ren
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07039__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _05265_ _05270_ _05291_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06406__X _01533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11363_ _05223_ _05224_ top.a1.dataIn\[19\] vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10075__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10594__A0 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13102_ clknet_leaf_116_clk _00666_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ net1955 net221 net398 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11294_ net892 top.a1.row1\[101\] _05168_ _01444_ vssd1 vssd1 vccd1 vccd1 _05169_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_210_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08988__B net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ clknet_leaf_3_clk _00597_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10245_ net2026 net221 net457 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1102 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09751__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ net233 net1571 net412 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_201_Left_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07762__A1 _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _04820_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_1
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__B2 top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload5_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ net1153 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_202_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12817_ clknet_leaf_3_clk _00381_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13797_ clknet_leaf_67_clk _01340_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07278__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ clknet_leaf_9_clk _00312_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09050__D _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_210_Left_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10821__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09019__A1 _03456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12679_ clknet_leaf_26_clk _00243_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13099__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold605 top.DUT.register\[25\]\[29\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 top.DUT.register\[6\]\[12\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 top.DUT.register\[13\]\[21\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 top.DUT.register\[15\]\[28\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold649 top.DUT.register\[9\]\[29\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ _01694_ net470 vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nand2_1
XANTENNA__10713__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ _04883_ _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07202__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__X _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ _01862_ _03922_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__nand2_1
XANTENNA__13593__Q top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06556__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08950__B1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ _01993_ net485 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07723_ top.DUT.register\[21\]\[1\] net575 net602 top.DUT.register\[10\]\[1\] _02849_
+ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__a221o_1
XANTENNA__06308__A2 _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout177_A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09522__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _02760_ _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__nand2_2
XFILLER_0_149_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06605_ net806 _01731_ _01624_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09258__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ _02691_ _02709_ net805 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_4
XFILLER_0_165_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1086_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09949__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _04370_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__or2_1
XANTENNA__07269__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06536_ net789 _01637_ _01643_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__and3_4
XANTENNA__07808__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _04302_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12375__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06467_ top.a1.instruction\[10\] top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ _01594_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _02879_ _03170_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06398_ _01496_ net793 _01503_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__and3_4
X_09186_ _04241_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08137_ net890 top.ru.state\[0\] net840 vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07441__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ net516 net289 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06795__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ top.DUT.register\[17\]\[11\] net646 net613 top.DUT.register\[14\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10623__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ net464 _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__nand2_8
XANTENNA__09194__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09733__A2 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06547__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _05834_ _05847_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a21oi_2
X_13720_ clknet_leaf_67_clk _00003_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_10932_ net154 net2246 net443 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07233__A _02339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13651_ clknet_leaf_83_clk _01210_ net1010 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10863_ net1656 net165 net352 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08048__B _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12602_ clknet_leaf_15_clk _00166_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ clknet_leaf_98_clk _01141_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10794_ net1678 net176 net445 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__mux2_1
X_12533_ clknet_leaf_90_clk _00097_ net998 vssd1 vssd1 vccd1 vccd1 top.pc\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12464_ clknet_leaf_97_clk top.ru.next_FetchedInstr\[16\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[16\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08064__A _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11415_ _05253_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2_1
X_12395_ clknet_leaf_84_clk _00031_ net1014 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07432__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ top.a1.dataIn\[27\] _05197_ top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 _05216_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__10533__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _05095_ _05115_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13016_ clknet_leaf_109_clk _00580_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10228_ net162 net2089 net405 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold2 _01179_ vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_146_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10159_ net166 net1925 net415 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07499__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08160__A1 _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13849_ net1114 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XANTENNA__06710__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09769__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ _02279_ _02404_ _02450_ _02496_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__or4b_1
XFILLER_0_18_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06321_ _01448_ _01330_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10708__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ net316 net285 _03296_ _04006_ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__o311a_1
X_06252_ net1324 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[28\] sky130_fd_sc_hd__and2_1
XFILLER_0_142_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07671__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06183_ top.a1.halfData\[2\] top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 _01412_
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_107_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold402 top.DUT.register\[30\]\[28\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 top.DUT.register\[30\]\[21\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 top.DUT.register\[24\]\[1\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 top.DUT.register\[17\]\[20\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__C1 _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 top.DUT.register\[14\]\[17\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 top.DUT.register\[16\]\[15\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 top.DUT.register\[24\]\[24\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net197 net1762 net436 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__mux2_1
XANTENNA__10443__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold479 top.DUT.register\[9\]\[16\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08421__B _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_2
Xfanout926 net933 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_55_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout937 net980 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_4
X_09873_ _04859_ _04862_ _04860_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__o21a_1
Xfanout948 net955 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_2
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08923__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net964 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_2
Xhold1102 top.DUT.register\[20\]\[7\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ _01865_ _03099_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_146_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 top.DUT.register\[10\]\[23\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1001_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 top.DUT.register\[8\]\[27\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 top.DUT.register\[6\]\[24\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 top.DUT.register\[19\]\[25\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net271 _03702_ _03858_ net273 _03855_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__o221a_1
Xhold1157 top.DUT.register\[20\]\[2\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_116_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1168 top.DUT.register\[4\]\[18\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__A1 top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1179 top.DUT.register\[18\]\[21\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _02206_ _02736_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__or2_1
XANTENNA__11286__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09252__B _04304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ net888 top.pc\[18\] net537 _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07637_ top.DUT.register\[8\]\[2\] net739 net700 top.DUT.register\[29\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout726_A _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06701__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ top.DUT.register\[11\]\[3\] net639 net548 top.DUT.register\[24\]\[3\] _02694_
+ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ top.pc\[15\] _04341_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__xnor2_1
X_06519_ _01644_ _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10618__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ top.DUT.register\[25\]\[5\] net624 net619 top.DUT.register\[26\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XANTENNA__08454__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__A1 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ net138 _04282_ _04291_ net911 vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__o211ai_1
XPHY_EDGE_ROW_125_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09169_ top.pc\[6\] _04210_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11200_ net1230 net530 _05087_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__a21o_1
XANTENNA__08171__X _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12180_ _01399_ _06046_ _06047_ _06048_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ net57 net858 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__and2_1
XANTENNA__10353__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 top.DUT.register\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 top.DUT.register\[18\]\[6\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net77 net864 net828 net1210 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__a22o_1
X_10013_ net229 net1586 net428 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_134_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10721__A0 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06940__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _05832_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__nand2_1
XANTENNA__08059__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13703_ clknet_leaf_73_clk _01251_ net1090 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ net210 net2136 net442 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11895_ net129 _05749_ _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13634_ clknet_leaf_61_clk net1242 net1101 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
X_10846_ net1378 net232 net350 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13565_ clknet_leaf_75_clk _01124_ net1088 vssd1 vssd1 vccd1 vccd1 top.a1.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_143_Left_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10777_ net2184 net245 net448 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__mux2_1
XANTENNA__10528__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12516_ clknet_leaf_70_clk _00008_ net1103 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13496_ clknet_leaf_111_clk _01060_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12447_ clknet_leaf_94_clk top.ru.next_FetchedData\[31\] net997 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07405__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12378_ net2351 net120 _00017_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
XANTENNA__06759__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ _05196_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__or2_1
XANTENNA__10263__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_Left_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06870_ top.DUT.register\[15\]\[22\] net707 net694 top.DUT.register\[21\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XANTENNA__08381__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06931__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08540_ net268 _03439_ _03443_ net272 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__B2 _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ net479 _03579_ _03586_ net520 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08684__A2 _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ top.DUT.register\[29\]\[6\] net703 net672 top.DUT.register\[16\]\[6\] _02547_
+ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07892__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_161_Left_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10946__B net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07353_ top.DUT.register\[29\]\[8\] net663 net627 top.DUT.register\[9\]\[8\] _02473_
+ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10438__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06304_ _01449_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XANTENNA__11123__A net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07284_ top.DUT.register\[20\]\[9\] net748 net726 top.DUT.register\[17\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06998__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09023_ _03727_ _04080_ _04082_ _04084_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__and4_1
X_06235_ net1252 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[11\] sky130_fd_sc_hd__and2_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1049_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_clk_X clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 top.DUT.register\[14\]\[10\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 top.lcd.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
Xhold232 top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 top.DUT.register\[19\]\[13\] vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 top.DUT.register\[14\]\[13\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold265 top.DUT.register\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 top.a1.data\[6\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 top.DUT.register\[28\]\[16\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09962__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 _01536_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
X_09925_ top.a1.instruction\[7\] top.a1.instruction\[8\] _04675_ vssd1 vssd1 vccd1
+ vccd1 _04916_ sky130_fd_sc_hd__nand3b_4
Xhold298 top.DUT.register\[30\]\[9\] vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout723 _01527_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
Xfanout734 _01522_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
Xfanout745 _01518_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout676_A _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 _01515_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_2
X_09856_ _04844_ _04847_ _04852_ _01586_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a31o_1
Xfanout767 net770 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10901__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 _01502_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 _01630_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_2
X_08807_ _01908_ net468 net487 vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__o21a_1
X_09787_ net834 _04402_ _04407_ net526 vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a2bb2o_1
X_06999_ top.DUT.register\[23\]\[11\] net698 net677 top.DUT.register\[18\]\[11\] _02125_
+ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06922__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ net478 _03836_ _03843_ net481 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12654__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _03034_ _03075_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10700_ net170 net1803 net378 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07883__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ _05506_ _05536_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_193_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10631_ net191 net2225 net392 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10348__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07635__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ clknet_leaf_23_clk _00914_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ net181 net2277 net357 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ top.lcd.cnt_500hz\[7\] _06106_ top.lcd.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1
+ _06108_ sky130_fd_sc_hd__a21o_1
XANTENNA__06989__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13281_ clknet_leaf_28_clk _00845_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12729__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ net208 net1567 net367 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__mux2_1
X_12232_ top.lcd.cnt_20ms\[5\] _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10083__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12163_ _06013_ _06018_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08061__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ net917 net1273 net855 _05043_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ _05959_ _05960_ _05954_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_207_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ net26 net842 net812 net2153 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_207_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08488__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06913__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11208__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ clknet_leaf_40_clk _00560_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12__f_clk_X clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11947_ _05784_ _05787_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07874__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _05707_ _05742_ _05710_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09112__S _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13617_ clknet_leaf_82_clk net1191 net1011 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
X_10829_ net2097 net170 net354 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__mux2_1
XANTENNA__10258__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07626__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ clknet_leaf_10_clk _01112_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13479_ clknet_leaf_8_clk _01043_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09348__A _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _01909_ _03097_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09710_ net836 _04269_ _04720_ top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _04724_
+ sky130_fd_sc_hd__a2bb2o_1
X_06922_ top.DUT.register\[8\]\[21\] net742 net694 top.DUT.register\[21\]\[21\] _02048_
+ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a221o_1
XANTENNA__10721__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _04657_ _04660_ _04666_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__or3_1
X_06853_ top.DUT.register\[14\]\[23\] net720 net685 top.DUT.register\[1\]\[23\] _01979_
+ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a221o_1
XANTENNA__06500__A top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06904__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__inv_2
X_06784_ top.DUT.register\[4\]\[24\] net769 _01539_ top.DUT.register\[13\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XANTENNA__09811__A top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ _03334_ _03619_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__a21o_1
XANTENNA__10379__D net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08657__A2 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ net2033 net840 net815 _03572_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07405_ top.DUT.register\[19\]\[7\] net631 net779 top.DUT.register\[15\]\[7\] _02522_
+ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_186_Right_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08385_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10168__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout424_A _04925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08146__B _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09957__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ top.DUT.register\[8\]\[8\] net739 _02451_ _02462_ vssd1 vssd1 vccd1 vccd1
+ _02463_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07267_ top.DUT.register\[4\]\[14\] net566 net558 top.DUT.register\[6\]\[14\] _02393_
+ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ _03678_ _03693_ _03698_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__nand3_1
X_06218_ top.Ren top.Wen vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__xnor2_1
X_07198_ top.DUT.register\[6\]\[15\] net764 net689 top.DUT.register\[3\]\[15\] _02322_
+ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_187_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08593__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout960_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net521 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06888__Y _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 _05078_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
Xfanout542 _01671_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10631__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _04011_ net343 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__nand2_1
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_8
Xfanout564 net567 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_4
Xfanout575 _01635_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_4
Xfanout586 _01512_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07506__A _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ net802 _04837_ _04838_ _04833_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a31o_1
Xfanout597 _01670_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ clknet_leaf_50_clk _00414_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11801_ _05610_ _05664_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_202_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12781_ clknet_leaf_32_clk _00345_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11732_ _05589_ _05600_ top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_138_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06409__X _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _05529_ _05531_ _05525_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a21o_1
XANTENNA__10078__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08056__B _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13402_ clknet_leaf_18_clk _00966_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10614_ net257 net1634 net389 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__mux2_1
X_11594_ _05441_ _05442_ _05416_ _05422_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ clknet_leaf_6_clk _00897_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10545_ top.DUT.register\[19\]\[31\] net140 net363 vssd1 vssd1 vccd1 vccd1 _00729_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10806__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ clknet_leaf_122_clk _00828_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10476_ net159 top.DUT.register\[17\]\[28\] net372 vssd1 vssd1 vccd1 vccd1 _00662_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08072__A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12215_ net1093 _04627_ net849 vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ clknet_leaf_30_clk _00759_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10915__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08584__A1 _02401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07387__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12146_ top.a1.dataIn\[2\] _06005_ _06012_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06595__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10541__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _05926_ _05929_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__or3_1
XANTENNA__08336__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__S _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output53_A net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ net7 net831 net830 net1707 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__a22o_1
XANTENNA__08887__A2 _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07770__A_N _02339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12979_ clknet_leaf_1_clk _00543_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07847__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07311__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08170_ _03295_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07121_ _02241_ _02243_ _02246_ _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_121_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13475__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07052_ top.DUT.register\[11\]\[10\] net755 net743 top.DUT.register\[31\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
XANTENNA__06822__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09521__A_N _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XANTENNA__10379__A_N net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06214__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13439__RESET_B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10451__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ _02909_ _03077_ _03074_ _03054_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_195_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08327__A1 _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06905_ top.DUT.register\[23\]\[22\] net562 net617 top.DUT.register\[30\]\[22\] _02016_
+ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_182_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07885_ _03002_ _03011_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout374_A _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ top.pad.keyCode\[0\] top.pad.keyCode\[2\] top.pad.keyCode\[3\] top.pad.keyCode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__or4b_1
X_06836_ top.DUT.register\[14\]\[23\] net611 net599 top.DUT.register\[10\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07550__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09555_ _04588_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nor2_1
XANTENNA__12378__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06767_ _01887_ _01889_ _01893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout541_A _01671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08506_ net281 _03580_ _03621_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07838__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09486_ top.pc\[25\] _04508_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__nor2_1
XANTENNA__08157__A _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06698_ top.DUT.register\[1\]\[26\] net687 net670 top.DUT.register\[5\]\[26\] _01824_
+ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a221o_1
XANTENNA__07302__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ _02496_ _03523_ _03548_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout806_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ _03486_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__nand2_2
XFILLER_0_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07319_ _02430_ _02432_ _02436_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__nor4_1
XFILLER_0_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10626__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08299_ net286 _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__or2_1
XANTENNA__09460__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10330_ net1466 net162 net397 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08015__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ net1523 net163 net454 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__mux2_1
X_12000_ _05842_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10192_ net169 net1864 net410 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10361__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 _04963_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_204_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 _04960_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_8
Xfanout372 _04958_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_4
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_8
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12902_ clknet_leaf_24_clk _00466_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13882_ net1132 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__08619__X _03731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07541__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ clknet_leaf_26_clk _00397_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ clknet_leaf_53_clk _00328_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08067__A _01929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__A2 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11715_ _05560_ _05584_ _05528_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12695_ clknet_leaf_106_clk _00259_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11646_ _05504_ _05508_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10536__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _05425_ _05433_ _05440_ _05442_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a22oi_1
Xclkbuf_leaf_103_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput36 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_13316_ clknet_leaf_39_clk _00880_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap506 net508 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10528_ net1870 net196 net363 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__mux2_1
Xhold809 top.DUT.register\[13\]\[13\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13247_ clknet_leaf_114_clk _00811_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08006__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ net219 net2142 net371 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
X_13178_ clknet_leaf_18_clk _00742_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10364__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06568__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10271__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _05994_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__nor2_1
XANTENNA__11864__A1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ top.DUT.register\[29\]\[0\] net663 net595 top.DUT.register\[27\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07532__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ top.DUT.register\[15\]\[28\] net706 net679 top.DUT.register\[13\]\[28\] _01747_
+ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06740__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09340_ _04385_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__or2_1
X_06552_ top.DUT.register\[6\]\[30\] net557 net604 top.DUT.register\[18\]\[30\] _01678_
+ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_47_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11115__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09271_ net138 _04312_ _04321_ _04322_ net911 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__o221a_1
X_06483_ _01607_ _01608_ net904 _01570_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_16_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08222_ net286 _03347_ _03292_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_16_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08264__X _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12414__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08153_ _03271_ _03278_ net308 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10446__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07599__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ _02225_ _02230_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__nor2_2
XANTENNA__08796__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08796__B2 _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _03207_ _03210_ net276 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ net809 net509 net463 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1031_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08440__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06512__X _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _04046_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nor2_1
XANTENNA__09970__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ top.DUT.register\[1\]\[16\] net656 net561 top.DUT.register\[23\]\[16\] _03063_
+ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a221o_1
XANTENNA__13202__RESET_B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A _01515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ top.DUT.register\[4\]\[17\] net767 net712 top.DUT.register\[30\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07523__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06819_ top.DUT.register\[2\]\[24\] net662 net554 top.DUT.register\[7\]\[24\] _01934_
+ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a221o_1
X_09607_ _04637_ _04638_ _04627_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ top.DUT.register\[4\]\[19\] net769 net669 top.DUT.register\[5\]\[19\] _02925_
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__a221o_1
XFILLER_0_210_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09538_ net133 _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _01929_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ _05316_ _05328_ _05341_ _05344_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4b_1
XFILLER_0_163_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12480_ clknet_leaf_95_clk top.ru.next_write_i net990 vssd1 vssd1 vccd1 vccd1 top.Wen
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08615__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _05298_ _05299_ _05294_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10356__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08787__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ _05205_ _05223_ _05224_ _05230_ _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06798__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ clknet_leaf_23_clk _00665_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ net2047 net225 net400 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ _05102_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13032_ clknet_leaf_35_clk _00596_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09736__B1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11138__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net1972 net223 net454 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
XANTENNA__06422__X _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1102 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10091__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ net235 top.DUT.register\[9\]\[8\] net409 vssd1 vssd1 vccd1 vccd1 _00386_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07762__A2 _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06970__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07253__X _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ net1152 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XANTENNA__12925__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06722__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11216__A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12816_ clknet_leaf_122_clk _00380_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13796_ clknet_leaf_65_clk _01339_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12747_ clknet_leaf_29_clk _00311_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09019__A2 _03537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12678_ clknet_leaf_19_clk _00242_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11629_ _05455_ _05456_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_42_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08778__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold606 top.DUT.register\[29\]\[3\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09059__C _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold617 top.DUT.register\[14\]\[31\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 top.DUT.register\[21\]\[28\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 top.DUT.register\[3\]\[31\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09727__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09356__A top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clk_X clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ net1453 net839 net815 _03940_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09075__B _03171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08771_ _03537_ _03542_ _03874_ net274 _03871_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o221a_2
XANTENNA__08950__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06961__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ top.DUT.register\[5\]\[1\] net547 net605 top.DUT.register\[18\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07505__A2 _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07653_ net495 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__inv_2
XFILLER_0_192_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06604_ _01726_ _01728_ _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__or3_4
X_07584_ _02690_ _02710_ net805 vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ top.pc\[15\] _04341_ top.pc\[16\] vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06535_ net789 _01634_ _01643_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_38_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11065__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout337_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1079_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ _04305_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06466_ top.a1.instruction\[29\] top.a1.instruction\[30\] top.a1.instruction\[31\]
+ _01566_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08205_ net474 vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08218__B1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13043__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ top.pc\[6\] _04210_ top.pc\[7\] vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10176__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06397_ top.DUT.register\[4\]\[30\] net770 net728 top.DUT.register\[10\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_190_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09965__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ net886 top.pc\[0\] _03261_ net539 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a22o_1
XANTENNA__09818__X _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08722__X _03829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _01929_ net294 vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__nand2_1
XANTENNA__10904__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ top.DUT.register\[29\]\[11\] net665 net658 top.DUT.register\[1\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a22o_1
XANTENNA__09718__B1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07057__Y _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07744__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net1389 net868 _02947_ net594 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _05825_ _05845_ _05834_ _05752_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_197_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10931_ net156 net1740 net443 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XANTENNA__06704__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13650_ clknet_leaf_84_clk _01209_ net1015 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
X_10862_ net1684 net168 net350 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12601_ clknet_leaf_36_clk _00165_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ clknet_leaf_98_clk _01140_ net981 vssd1 vssd1 vccd1 vccd1 top.ramload\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10793_ top.DUT.register\[27\]\[22\] net185 net448 vssd1 vssd1 vccd1 vccd1 _00976_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ clknet_leaf_88_clk _00096_ net1005 vssd1 vssd1 vccd1 vccd1 top.pc\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08345__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10086__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ clknet_leaf_100_clk top.ru.next_FetchedInstr\[15\] net997 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _05248_ _05256_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and2_1
X_12394_ clknet_leaf_88_clk _00030_ net1005 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08632__X _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11345_ _05212_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10814__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07983__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09176__A _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ top.lcd.nextState\[4\] net882 net879 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o21ba_1
X_13015_ clknet_leaf_17_clk _00579_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10227_ net164 net1807 net407 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ net170 net1832 net416 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 top.pad.button_control.debounce vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06943__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10089_ net171 net2295 net418 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13848_ net1113 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08448__B1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ clknet_leaf_64_clk _01322_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09645__C1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06320_ _01459_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07120__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08255__A _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06251_ net1325 net872 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[27\] sky130_fd_sc_hd__and2_1
XFILLER_0_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06182_ net893 _00017_ _01409_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold403 top.DUT.register\[28\]\[19\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 top.DUT.register\[7\]\[27\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10724__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold425 top.DUT.register\[16\]\[29\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08261__Y _03386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold436 top.DUT.register\[6\]\[16\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold447 top.DUT.register\[18\]\[13\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 top.DUT.register\[30\]\[3\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ net201 net1964 net435 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__mux2_1
Xhold469 top.DUT.register\[8\]\[10\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout905 top.a1.instruction\[4\] vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
Xfanout916 net918 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_2
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
X_09872_ net167 net2118 net440 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07187__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
Xfanout949 net955 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
Xhold1103 top.DUT.register\[26\]\[2\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_146_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 top.DUT.register\[6\]\[8\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1125 top.DUT.register\[20\]\[27\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 top.DUT.register\[25\]\[18\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__inv_2
Xhold1147 top.lcd.currentState\[5\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 top.DUT.register\[30\]\[29\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 top.DUT.register\[8\]\[30\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ top.a1.instruction\[22\] _02208_ net529 vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__o21a_1
XANTENNA__08687__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ net471 _03784_ _03793_ _03783_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_179_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08149__B _03012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_A _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10494__A0 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ top.DUT.register\[12\]\[2\] net580 net667 top.DUT.register\[5\]\[2\] _02762_
+ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ top.DUT.register\[9\]\[3\] net627 net611 top.DUT.register\[14\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09306_ top.i_ready top.pc\[14\] _04355_ net899 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__o211a_1
X_06518_ top.a1.instruction\[20\] top.a1.instruction\[21\] net900 _01626_ vssd1 vssd1
+ vccd1 vccd1 _01645_ sky130_fd_sc_hd__o31a_1
XFILLER_0_63_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07498_ top.DUT.register\[19\]\[5\] net631 net781 top.DUT.register\[31\]\[5\] _02624_
+ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a221o_1
XANTENNA__07111__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ net134 _04285_ _04290_ net819 vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__o22a_1
XANTENNA__13635__RESET_B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06449_ top.a1.instruction\[12\] net902 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_157_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09695__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ net908 top.pc\[5\] _04226_ net898 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08119_ _02184_ net295 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__nand2_1
XANTENNA__10634__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ _04159_ _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_170_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ net914 net1299 net854 _05051_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a31o_1
Xhold970 top.DUT.register\[25\]\[1\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 top.ramaddr\[27\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold992 top.DUT.register\[23\]\[30\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ net76 net864 net828 net1161 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a22o_1
XANTENNA__07178__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ net181 net1619 net425 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XANTENNA__07717__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06925__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _05798_ _05822_ _05823_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13702_ clknet_leaf_73_clk _01250_ net1093 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ net219 net2099 net443 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
X_11894_ _05730_ _05733_ _05727_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07350__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10845_ net1624 net237 net349 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
X_13633_ clknet_leaf_98_clk net1259 net981 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10809__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10776_ net2071 net248 net445 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__mux2_1
X_13564_ clknet_leaf_75_clk _01123_ net1088 vssd1 vssd1 vccd1 vccd1 top.a1.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06345__C_N net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12515_ clknet_leaf_45_clk _00082_ net1081 vssd1 vssd1 vccd1 vccd1 top.ramstore\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11213__B top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ clknet_leaf_77_clk _01059_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ clknet_leaf_95_clk top.ru.next_FetchedData\[30\] net991 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[30\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__08362__X _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12377_ top.pad.keyCode\[6\] net119 _00017_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10544__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11328_ _05194_ _05195_ top.a1.dataIn\[26\] vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10960__B2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11259_ net1266 net824 _05137_ net1090 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__o211a_1
XANTENNA__07169__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06916__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_74_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_187_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08470_ _02450_ net470 _03584_ net522 _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_141_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06993__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ top.DUT.register\[19\]\[6\] net733 net715 top.DUT.register\[30\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06695__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07352_ top.DUT.register\[8\]\[8\] net568 net552 top.DUT.register\[7\]\[8\] _02478_
+ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_174_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06303_ net2307 _01445_ _01446_ top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 _01449_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07283_ top.DUT.register\[30\]\[9\] net713 net686 top.DUT.register\[1\]\[9\] _02409_
+ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a221o_1
XANTENNA__06217__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ net273 _03426_ _03565_ net317 _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__o221a_1
X_06234_ net2111 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[10\] sky130_fd_sc_hd__and2_1
XFILLER_0_143_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold200 net88 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10454__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06165_ top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold211 top.DUT.register\[13\]\[19\] vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 top.DUT.register\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold233 top.DUT.register\[12\]\[10\] vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 top.DUT.register\[23\]\[15\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold266 top.DUT.register\[23\]\[18\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 top.DUT.register\[13\]\[7\] vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09149__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold288 top.DUT.register\[19\]\[22\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 top.DUT.register\[13\]\[5\] vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout702 _01536_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_8
X_09924_ net141 net1904 net439 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__mux2_1
Xfanout713 _01531_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_4
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout724 _01525_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_8
Xfanout735 _01521_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
Xfanout746 _01518_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_2
XANTENNA__09544__A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06520__X _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _04844_ _04847_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a21oi_1
Xfanout757 _01515_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06907__B1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 net780 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_4
XANTENNA_fanout669_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net481 _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__or2_1
XANTENNA__09263__B _04304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06998_ top.DUT.register\[22\]\[11\] net753 net707 top.DUT.register\[15\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a22o_1
X_09786_ _04776_ _04780_ _04789_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__or3b_1
XANTENNA__07580__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ _03478_ _03542_ _03841_ net274 _03842_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__o221a_1
XANTENNA__11259__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ net1328 net840 net815 _03777_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07332__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13381__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12208__A1 top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ top.DUT.register\[28\]\[2\] net651 net540 top.DUT.register\[22\]\[2\] _02740_
+ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a221o_1
XANTENNA__06686__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10629__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ net473 _03692_ _03711_ net476 _03706_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ net206 net1592 net391 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ net197 net2314 net358 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ top.lcd.cnt_500hz\[7\] _06106_ _06107_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__o21a_1
XANTENNA__09278__X _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ clknet_leaf_44_clk _00844_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ net222 net2087 net368 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12231_ top.lcd.cnt_20ms\[4\] top.lcd.cnt_20ms\[3\] _06063_ vssd1 vssd1 vccd1 vccd1
+ _06064_ sky130_fd_sc_hd__and3_1
XANTENNA__09388__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12162_ top.a1.dataIn\[2\] _06011_ _06012_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__o21ba_1
X_11113_ net47 net857 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__and2_1
XANTENNA__06610__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ _05959_ _05960_ _05952_ _05953_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ net25 net831 _05024_ net1362 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__a22o_1
XANTENNA__09454__A _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08363__A2 _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07571__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12995_ clknet_leaf_33_clk _00559_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09312__A1 _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11946_ _05776_ _05782_ _05786_ _05790_ _05777_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a41o_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06677__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10539__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ _05736_ _05741_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__a21o_1
X_13616_ clknet_leaf_98_clk net1184 net981 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828_ net1410 net172 net355 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__mux2_1
XANTENNA__06318__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06429__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ clknet_leaf_30_clk _01111_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10759_ net193 top.DUT.register\[26\]\[20\] net376 vssd1 vssd1 vccd1 vccd1 _00942_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13478_ clknet_leaf_9_clk _01042_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12429_ clknet_leaf_96_clk top.ru.next_FetchedData\[13\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[13\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09348__B _03011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07929__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07149__A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ _01930_ _01949_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06601__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06921_ top.DUT.register\[22\]\[21\] net753 net710 top.DUT.register\[9\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__09551__A1 top.a1.instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ _04643_ _04653_ _04646_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a21oi_1
X_06852_ top.DUT.register\[25\]\[23\] net771 net731 top.DUT.register\[19\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a22o_1
X_09571_ top.a1.instruction\[30\] net822 _04424_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__o21a_2
X_06783_ top.DUT.register\[26\]\[24\] net761 net749 top.DUT.register\[20\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_47_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08522_ _03635_ _03637_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11110__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07314__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08965__A1_N net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ net887 top.pc\[8\] net536 _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a22o_1
XANTENNA__06668__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07404_ top.DUT.register\[8\]\[7\] net568 net607 top.DUT.register\[12\]\[7\] _02530_
+ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ _03454_ _03504_ net278 vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07335_ top.DUT.register\[28\]\[8\] net584 net667 top.DUT.register\[5\]\[8\] _02461_
+ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1061_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout417_A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07093__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ top.DUT.register\[21\]\[14\] net575 net634 top.DUT.register\[19\]\[14\] _02392_
+ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a221o_1
XANTENNA__06515__X _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09005_ _03254_ _03351_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06217_ net1 net855 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10184__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06840__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07197_ top.DUT.register\[30\]\[15\] net713 net701 top.DUT.register\[29\]\[15\] _02323_
+ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a221o_1
XANTENNA__09973__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_203_Right_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout521 _03258_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
Xfanout532 _05064_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
X_09907_ net152 net1957 net439 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__mux2_1
Xfanout543 _01671_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_4
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net566 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10688__A0 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 _01633_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_8
Xfanout587 _01512_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
X_09838_ _04821_ _04826_ _04836_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__nand3_1
Xfanout598 _01670_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07553__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ net227 net2215 net437 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11800_ _05663_ _05666_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__or3b_1
XFILLER_0_197_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ clknet_leaf_10_clk _00344_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07305__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _05589_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nand2_1
XANTENNA__06659__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11662_ _05529_ _05531_ _05525_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13401_ clknet_leaf_37_clk _00965_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ net261 net2037 net389 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__mux2_1
XANTENNA__11979__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07608__B2 top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _05441_ _05442_ _05416_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13332_ clknet_leaf_46_clk _00896_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10544_ net2191 net146 net362 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__mux2_1
XANTENNA__10094__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06831__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ net163 top.DUT.register\[17\]\[27\] net369 vssd1 vssd1 vccd1 vccd1 _00661_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13277__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13263_ clknet_leaf_21_clk _00827_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12214_ net1316 net846 net814 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__a21o_1
X_13194_ clknet_leaf_40_clk _00758_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08584__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__A1 top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ _05992_ _06002_ _05990_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__a21o_1
XANTENNA__10822__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07792__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _05937_ _05941_ _05942_ _05943_ _05935_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__o41a_2
XANTENNA__08336__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ net6 net841 net811 net1320 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__o22a_1
XANTENNA__07544__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07703__Y _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12978_ clknet_leaf_50_clk _00542_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10269__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _05770_ _05791_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13859__1150 vssd1 vssd1 vccd1 vccd1 net1150 _13859__1150/LO sky130_fd_sc_hd__conb_1
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07120_ top.DUT.register\[19\]\[12\] net732 net718 top.DUT.register\[2\]\[12\] _02244_
+ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09359__A top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07051_ top.DUT.register\[28\]\[10\] net584 _02168_ _02177_ vssd1 vssd1 vccd1 vccd1
+ _02178_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_136_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06822__A2 _01948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_88_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_113_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10732__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _02928_ _02948_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_182_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06904_ top.DUT.register\[28\]\[22\] net654 net570 top.DUT.register\[8\]\[22\] _02030_
+ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_182_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07884_ _03003_ _03006_ _03008_ _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__or4_4
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _04647_ _04651_ _01472_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_207_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06889__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06835_ top.DUT.register\[4\]\[23\] net564 net619 top.DUT.register\[26\]\[23\] _01961_
+ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout367_A _04959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09554_ _01713_ _04587_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and2b_1
X_06766_ top.DUT.register\[21\]\[25\] net575 _01890_ _01892_ vssd1 vssd1 vccd1 vccd1
+ _01893_ sky130_fd_sc_hd__a211o_1
XFILLER_0_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08505_ net288 _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06697_ top.DUT.register\[14\]\[26\] net722 net673 top.DUT.register\[16\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a22o_1
X_09485_ _01587_ _04523_ _04178_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout534_A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__SET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ _03523_ _03548_ _02496_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08367_ net473 _03465_ _03488_ net476 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07318_ _02438_ _02440_ _02442_ _02444_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__or4_1
XFILLER_0_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08263__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _03313_ _03317_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07249_ top.DUT.register\[22\]\[14\] net754 net679 top.DUT.register\[13\]\[14\] _02366_
+ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a221o_1
XANTENNA__06813__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10260_ net1520 net164 net457 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ net173 net1929 net410 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XANTENNA__10642__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
Xfanout351 _04963_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_204_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout362 _04960_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_2
Xfanout373 _04952_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_8
Xfanout384 _04947_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07526__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_6
X_12901_ clknet_leaf_117_clk _00465_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13881_ net1131 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_107_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ clknet_leaf_44_clk _00396_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13149__RESET_B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12763_ clknet_leaf_57_clk _00327_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10089__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11714_ top.a1.dataIn\[8\] _05582_ _05583_ top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1
+ _05584_ sky130_fd_sc_hd__or4b_1
XFILLER_0_194_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12694_ clknet_leaf_119_clk _00258_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11645_ _05510_ _05511_ _05513_ _05466_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__o211ai_2
XANTENNA__10817__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11576_ _05444_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or2_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
X_13315_ clknet_leaf_41_clk _00879_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11221__B top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_2
X_10527_ net1403 net199 net363 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10458_ net224 net1613 net370 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
X_13246_ clknet_leaf_14_clk _00810_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08811__A _01909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10552__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ clknet_leaf_36_clk _00741_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10389_ net240 net1891 net327 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ _05987_ net126 _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12059_ _05911_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06620_ top.DUT.register\[31\]\[28\] net746 net670 top.DUT.register\[5\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a22o_1
XANTENNA__11236__X _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13501__RESET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08258__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06551_ top.DUT.register\[11\]\[30\] net640 net549 top.DUT.register\[24\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09270_ _04319_ _04320_ _01618_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06482_ top.a1.instruction\[5\] _01570_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__nor2_1
XANTENNA__08493__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08221_ net293 net490 vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10727__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08152_ _03274_ _03277_ net282 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07103_ _02214_ _02226_ _02227_ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08083_ _03208_ _03209_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__nand2_1
XANTENNA__08796__A2 top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07034_ _02147_ _02158_ _02159_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__nor4_1
XFILLER_0_113_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10462__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1024_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ net895 _02835_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_149_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ top.DUT.register\[18\]\[16\] net604 net595 top.DUT.register\[27\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ top.DUT.register\[8\]\[17\] net739 net704 top.DUT.register\[15\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout749_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ top.a1.state\[2\] top.a1.state\[1\] net893 _04629_ vssd1 vssd1 vccd1 vccd1
+ _04638_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06818_ top.DUT.register\[9\]\[24\] net628 net547 top.DUT.register\[5\]\[24\] _01944_
+ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a221o_1
X_07798_ top.DUT.register\[11\]\[19\] net757 net724 top.DUT.register\[17\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09537_ _04569_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__xor2_1
X_06749_ top.DUT.register\[11\]\[25\] net756 net695 top.DUT.register\[21\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ top.a1.instruction\[24\] net821 _04424_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__o21a_2
XANTENNA__07287__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08419_ _03177_ _03524_ _03523_ net483 vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10637__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ net821 _02186_ _04424_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__o21a_2
X_11430_ _05298_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__nand2_1
XANTENNA__07039__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ top.a1.dataIn\[21\] _05210_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ clknet_leaf_8_clk _00664_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10312_ net1481 net232 net400 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
XANTENNA__07995__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11292_ net879 net881 top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08631__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10243_ net1365 net232 net455 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
X_13031_ clknet_leaf_7_clk _00595_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09736__B2 top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A1 top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1109 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
X_10174_ net242 net1308 net412 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
Xfanout170 _04858_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_2
Xfanout181 net182 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout192 _04811_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09462__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13864_ net1125 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XANTENNA__08078__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11216__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12815_ clknet_leaf_21_clk _00379_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ clknet_leaf_66_clk _01338_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12746_ clknet_leaf_37_clk _00310_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07278__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__B2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08806__A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10547__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ clknet_leaf_120_clk _00241_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11628_ _05451_ _05496_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_42_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08778__A2 _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11559_ _05368_ _05427_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09059__D net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 top.DUT.register\[8\]\[31\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07986__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold618 top.DUT.register\[17\]\[0\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 top.DUT.register\[31\]\[27\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07450__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09727__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10282__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ clknet_leaf_33_clk _00793_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07738__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07202__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08950__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ _03801_ _03873_ net307 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__mux2_1
XANTENNA__09372__A top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _02839_ _02841_ _02843_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__or4_1
XANTENNA__08702__A2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _02770_ _02771_ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__nor3_1
XANTENNA__07910__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06603_ top.DUT.register\[5\]\[29\] net546 net597 top.DUT.register\[27\]\[29\] _01729_
+ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a221o_1
X_07583_ _02709_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__inv_2
X_06534_ _01632_ _01644_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_4
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09322_ top.pc\[15\] top.pc\[16\] _04341_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__and3_1
XANTENNA__07269__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06465_ _01590_ _01591_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__and2_1
X_09253_ _02142_ _04304_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__and2_1
XANTENNA__10457__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout232_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12982__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ _03165_ _03173_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nand2_1
XANTENNA__08218__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09184_ top.pc\[6\] top.pc\[7\] _04210_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__and3_1
X_06396_ _01498_ _01499_ net790 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__and3_2
XFILLER_0_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ top.ru.next_write_i _00005_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08066_ _03191_ _03192_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__nand2_1
XANTENNA__07441__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06523__X _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ top.DUT.register\[3\]\[11\] net787 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout699_A _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__B2 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09981__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06401__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _02989_ net591 net1239 net869 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__a2bb2o_1
X_07919_ top.DUT.register\[10\]\[16\] net728 net686 top.DUT.register\[1\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ net1331 net839 net817 _03996_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_197_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ net161 net1789 net441 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07901__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10861_ net1920 net171 net349 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12600_ clknet_leaf_108_clk _00164_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07801__Y _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13580_ clknet_leaf_98_clk _01139_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10792_ net1364 net188 net447 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12531_ clknet_leaf_88_clk _00095_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[14\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__10367__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12462_ clknet_leaf_97_clk top.ru.next_FetchedInstr\[14\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11413_ _05246_ _05280_ _05281_ _05279_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__nor4b_1
X_12393_ clknet_leaf_82_clk _00029_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07432__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _05200_ _05213_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__or2_2
XANTENNA__08361__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09176__B _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ top.a1.row2\[35\] _05107_ _05119_ top.a1.row1\[19\] _05151_ vssd1 vssd1 vccd1
+ vccd1 _05152_ sky130_fd_sc_hd__a221o_1
X_13014_ clknet_leaf_2_clk _00578_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10226_ net168 net2055 net406 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__mux2_1
XANTENNA__10830__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ net171 net1721 net416 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 top.busy_o vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09192__A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ net177 net2091 net417 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XANTENNA__07499__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ net1112 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_202_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08448__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13778_ clknet_leaf_64_clk net1250 vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07440__A _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12729_ clknet_leaf_37_clk _00293_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10277__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06250_ net1675 net873 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[26\] sky130_fd_sc_hd__and2_1
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07671__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06181_ net893 _01409_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__and2_2
XFILLER_0_20_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold404 top.DUT.register\[6\]\[10\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold415 top.DUT.register\[27\]\[11\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08620__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 top.DUT.register\[4\]\[16\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08620__B2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10963__C1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold437 top.DUT.register\[8\]\[13\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 top.DUT.register\[6\]\[29\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06631__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold459 top.DUT.register\[4\]\[15\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ net210 net2054 net434 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout917 net918 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_2
X_09871_ _03937_ net341 net337 _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__o211a_4
XFILLER_0_110_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout928 net933 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09581__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _01865_ _03921_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__or2_1
XANTENNA__10740__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 top.DUT.register\[16\]\[12\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 top.DUT.register\[18\]\[24\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 top.DUT.register\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 top.DUT.register\[30\]\[0\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ _03787_ _03857_ net304 vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__mux2_1
Xhold1148 top.DUT.register\[4\]\[20\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout182_A _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__B1 _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 top.DUT.register\[28\]\[4\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07704_ net291 net467 vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__nand2_1
X_08684_ net522 _03790_ _03792_ _03785_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_205_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06698__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ top.DUT.register\[6\]\[2\] net763 net708 top.DUT.register\[9\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08439__B2 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07566_ top.DUT.register\[27\]\[3\] net595 net540 top.DUT.register\[22\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_192_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09305_ net138 _04343_ _04354_ net911 vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_158_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06517_ _01643_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10187__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07497_ top.DUT.register\[3\]\[5\] net785 net779 top.DUT.register\[15\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout614_A _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__X _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ _04288_ _04289_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06448_ top.a1.instruction\[25\] top.a1.instruction\[26\] _01574_ vssd1 vssd1 vccd1
+ vccd1 _01575_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06870__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06379_ top.a1.instruction\[18\] net810 top.a1.instruction\[17\] vssd1 vssd1 vccd1
+ vccd1 _01506_ sky130_fd_sc_hd__and3b_2
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ net137 _04212_ _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10915__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08452__Y _03571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08118_ _03241_ _03244_ net279 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13675__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _02739_ _02780_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_170_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ _03171_ _03173_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__and3_1
Xhold960 wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 top.DUT.register\[23\]\[23\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net75 net862 net826 net1206 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a22o_1
Xhold982 top.DUT.register\[17\]\[11\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold993 top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__D1 _03343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ net195 net1913 net426 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
XANTENNA__08914__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10650__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08127__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11962_ _05822_ _05823_ _05798_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_86_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ clknet_leaf_72_clk _01249_ net1096 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[109\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ net224 net1851 net441 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06689__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11893_ _05761_ _05762_ _05760_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__mux2_1
XANTENNA__12557__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13632_ clknet_leaf_61_clk net1189 net1100 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10844_ net1702 net241 net350 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13563_ clknet_leaf_75_clk _01122_ net1090 vssd1 vssd1 vccd1 vccd1 top.a1.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10775_ net1921 net253 net447 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12514_ clknet_leaf_45_clk _00081_ net1081 vssd1 vssd1 vccd1 vccd1 top.ramstore\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11213__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ clknet_leaf_2_clk _01058_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06861__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12445_ clknet_leaf_95_clk top.ru.next_FetchedData\[29\] net991 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[29\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10825__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07405__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ net2292 net118 _00017_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06613__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ top.a1.dataIn\[26\] _05194_ _05195_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09915__A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11258_ _05131_ _05133_ _05135_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12162__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ net237 net1748 net405 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__mux2_1
XANTENNA__10560__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net850 _05068_ net531 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__and3_1
XFILLER_0_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10132__Y _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12980__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08537__Y _03652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ top.DUT.register\[11\]\[6\] net758 net737 top.DUT.register\[24\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XANTENNA__07892__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11425__B1 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ top.DUT.register\[1\]\[8\] net655 net623 top.DUT.register\[25\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06302_ _01448_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ top.DUT.register\[6\]\[9\] net764 net716 top.DUT.register\[2\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_75_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09021_ net273 _03386_ _03190_ _03183_ _03343_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__o2111a_1
X_06233_ net1302 net871 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[9\] sky130_fd_sc_hd__and2_1
XANTENNA__06852__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06164_ top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XANTENNA__09097__A _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 _01190_ vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 top.DUT.register\[11\]\[15\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold223 top.DUT.register\[12\]\[15\] vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 top.DUT.register\[25\]\[15\] vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 top.DUT.register\[28\]\[21\] vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold256 top.DUT.register\[23\]\[10\] vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 top.DUT.register\[27\]\[12\] vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 top.DUT.register\[31\]\[1\] vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _04028_ net342 net339 _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__o211a_2
Xfanout703 _01536_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold289 top.DUT.register\[27\]\[3\] vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout714 _01531_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
Xfanout725 _01525_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 _01521_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10470__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ top.pc\[25\] _04518_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__xnor2_1
Xfanout747 _01517_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_8
Xfanout758 _01515_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_84_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06907__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ _03583_ _03906_ net322 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XANTENNA__12959__Q top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07345__A _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09785_ _04776_ _04780_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__o21bai_1
X_06997_ top.DUT.register\[27\]\[11\] net778 net762 top.DUT.register\[26\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout564_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09306__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08736_ net271 _03681_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13526__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_A _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ net890 top.pc\[17\] net539 _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07618_ top.DUT.register\[23\]\[2\] net560 net544 top.DUT.register\[5\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__A _02380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07883__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08598_ _03709_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11314__B top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ top.DUT.register\[18\]\[4\] net676 _02671_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _02676_ sky130_fd_sc_hd__a211o_1
XANTENNA__09085__B2 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07096__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07635__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ net199 net1795 net358 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__mux2_1
XANTENNA__06843__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _04270_ _04273_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_20_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10645__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10491_ net225 net2115 net366 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ top.lcd.cnt_20ms\[2\] top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] vssd1 vssd1
+ vccd1 vccd1 _06063_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ net125 _06030_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_112_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ net917 net1786 net852 _05042_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a31o_1
XANTENNA__09735__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12092_ _05959_ _05960_ _05952_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21o_1
Xhold790 top.DUT.register\[31\]\[20\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ net23 net842 net812 net1363 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_207_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07020__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12994_ clknet_leaf_42_clk _00558_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ _05797_ _05798_ _05799_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__a31o_1
XFILLER_0_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _05743_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__nand2_1
XANTENNA__07874__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13615_ clknet_leaf_98_clk net1268 net982 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
X_10827_ net1512 net177 net353 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07087__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13546_ clknet_leaf_34_clk _01110_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07626__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10758_ net203 net2218 net375 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__A _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06834__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13477_ clknet_leaf_116_clk _01041_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13526__RESET_B net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ net196 net1503 net379 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
X_12428_ clknet_leaf_95_clk top.ru.next_FetchedData\[12\] net990 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11186__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ net1348 _06142_ net795 vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07149__B _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06920_ top.DUT.register\[17\]\[21\] net724 net677 top.DUT.register\[18\]\[21\] _02046_
+ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a221o_1
XANTENNA__10290__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10146__A0 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07011__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13549__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ top.DUT.register\[11\]\[23\] net755 net667 top.DUT.register\[5\]\[23\] _01977_
+ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a221o_1
XANTENNA__09083__C _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06365__A2 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09570_ _04602_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__nand2b_1
X_06782_ _01907_ _01908_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nor2_2
X_08521_ net480 _03630_ _03634_ net477 _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07171__Y _02298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ _03569_ _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__nand2_2
XFILLER_0_148_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07403_ top.DUT.register\[24\]\[7\] net549 net596 top.DUT.register\[27\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08383_ _03227_ _03231_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout145_A _04908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ top.DUT.register\[20\]\[8\] net747 net708 top.DUT.register\[9\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07617__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10973__B net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10465__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07265_ top.DUT.register\[3\]\[14\] net788 _02391_ vssd1 vssd1 vccd1 vccd1 _02392_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout312_A _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _03596_ _04065_ _03753_ _03575_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__or4b_1
XFILLER_0_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06216_ wb.curr_state\[1\] wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__or2_1
X_07196_ top.DUT.register\[4\]\[15\] net767 net693 top.DUT.register\[21\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07250__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout681_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ _03994_ net344 _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a21oi_4
Xfanout522 _03183_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout533 _05064_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_2
Xfanout544 _01665_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_8
Xfanout555 _01654_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_4
XANTENNA__07002__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_8
X_09837_ _04821_ _04826_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a21o_1
Xfanout577 _01633_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
Xfanout588 _06098_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 _01669_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout946_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12916__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _03757_ net342 net339 _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__o211a_2
XFILLER_0_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08719_ _03456_ _03542_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_202_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _03552_ net340 net336 _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11730_ _05595_ _05597_ _05588_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a21o_2
XFILLER_0_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07856__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08775__B1_N _03878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ _05487_ _05526_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ clknet_leaf_110_clk _00964_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net263 net1659 net391 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__mux2_1
X_11592_ _05432_ _05454_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08634__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ clknet_leaf_5_clk _00895_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ net1871 net152 net363 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13262_ clknet_leaf_116_clk _00826_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10474_ net164 net2139 net371 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12213_ net2347 net849 _04976_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ clknet_leaf_12_clk _00757_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12144_ top.a1.dataIn\[2\] _06012_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07241__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06595__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12075_ _05941_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__or2_1
XANTENNA__08336__A3 _03456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ net5 net842 net812 net1287 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__o22a_1
XANTENNA__11219__B top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12596__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12977_ clknet_leaf_110_clk _00541_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11928_ _05729_ _05751_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07847__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ top.a1.dataIn\[6\] _05713_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06807__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13529_ clknet_leaf_36_clk _01093_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10285__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07050_ top.DUT.register\[29\]\[10\] net700 net692 top.DUT.register\[21\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_149_Left_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_121_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08980__B1 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__B _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _03012_ _03032_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__nand2b_1
X_06903_ top.DUT.register\[21\]\[22\] net574 net553 top.DUT.register\[7\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_182_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11129__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07883_ top.DUT.register\[17\]\[17\] net726 net716 top.DUT.register\[2\]\[17\] _03009_
+ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07535__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__B1 _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ top.pad.keyCode\[5\] top.pad.keyCode\[4\] top.pad.keyCode\[6\] top.pad.keyCode\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__or4b_2
X_06834_ top.DUT.register\[20\]\[23\] net576 net572 top.DUT.register\[21\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_158_Left_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08719__A _03456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__B net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _04587_ _01713_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__and2b_1
XANTENNA__08256__A2_N _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06765_ top.DUT.register\[2\]\[25\] net662 net569 top.DUT.register\[8\]\[25\] _01891_
+ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout262_A _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__B2 _01588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08504_ _03304_ _03308_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07838__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _04521_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06696_ top.DUT.register\[26\]\[26\] net762 net682 top.DUT.register\[7\]\[26\] _01822_
+ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ _02496_ _02893_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__xor2_1
XFILLER_0_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08366_ _02636_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__xor2_1
XANTENNA__06526__X _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07317_ top.DUT.register\[4\]\[9\] net567 net545 top.DUT.register\[5\]\[9\] _02443_
+ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10195__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ _03419_ _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__nand2_1
XANTENNA__08173__B _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07471__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07248_ top.DUT.register\[18\]\[14\] net676 net669 top.DUT.register\[5\]\[14\] _02374_
+ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout896_A top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09740__A1_N net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09212__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08015__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ top.DUT.register\[20\]\[13\] net578 _02303_ _02305_ vssd1 vssd1 vccd1 vccd1
+ _02306_ sky130_fd_sc_hd__a211o_1
X_10190_ net176 net1729 net409 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07517__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 _04956_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_8
Xfanout341 net342 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout352 _04963_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_204_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout363 _04960_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_8
Xfanout374 _04952_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_4
Xfanout385 _04945_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_8
X_12900_ clknet_leaf_39_clk _00464_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout396 _04943_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_4
X_13880_ top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09732__B _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ clknet_leaf_115_clk _00395_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12762_ clknet_leaf_16_clk _00326_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07829__A2 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07820__X _02947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11713_ top.a1.dataIn\[7\] top.a1.dataIn\[6\] top.a1.dataIn\[5\] top.a1.dataIn\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_120_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12693_ clknet_leaf_6_clk _00257_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11644_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__inv_2
XFILLER_0_204_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11575_ top.a1.dataIn\[13\] _05441_ _05442_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__and3_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A1 _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
X_13314_ clknet_leaf_43_clk _00878_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput38 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
X_10526_ net2158 net207 net362 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13245_ clknet_leaf_112_clk _00809_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10457_ net233 net2177 net370 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
XANTENNA__08006__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10833__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07214__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ clknet_leaf_109_clk _00740_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10388_ net243 net1916 net329 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07765__A1 _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06568__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _05979_ _05995_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12058_ _05923_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nand2_2
XANTENNA__08714__B1 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net1251 _05021_ net535 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__mux2_1
XANTENNA__08539__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06740__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06550_ top.DUT.register\[20\]\[30\] net577 net630 top.DUT.register\[9\]\[30\] _01676_
+ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06481_ _01387_ _01480_ _01577_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08493__A2 _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08220_ net473 _03336_ _03345_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_138_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _03275_ _03276_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07102_ top.DUT.register\[21\]\[10\] net572 net615 top.DUT.register\[30\]\[10\] _02228_
+ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08082_ _02056_ net294 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07033_ top.DUT.register\[4\]\[11\] net565 net625 top.DUT.register\[25\]\[11\] _02149_
+ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a221o_1
XANTENNA__10743__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07205__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__B1 _02709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ net895 _02835_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1017_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13117__CLK clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ top.DUT.register\[21\]\[16\] net573 net635 top.DUT.register\[16\]\[16\] _03061_
+ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_149_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07866_ _02991_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__nor2_2
X_09605_ _04631_ _04633_ _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_162_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06817_ top.DUT.register\[29\]\[24\] net664 net549 top.DUT.register\[24\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout644_A _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07797_ top.DUT.register\[15\]\[19\] net706 _02910_ _02923_ vssd1 vssd1 vccd1 vccd1
+ _02924_ sky130_fd_sc_hd__a211o_1
XANTENNA__09979__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _04570_ _04571_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nand2b_1
X_06748_ _01871_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ net136 _04506_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08484__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06679_ top.DUT.register\[23\]\[27\] net560 net608 top.DUT.register\[12\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__a22o_1
XANTENNA__10918__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08418_ _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__inv_2
XANTENNA__06495__A1 top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13211__RESET_B net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ _04438_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ net308 _03278_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07444__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ _05205_ _05210_ _05223_ _05224_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_132_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06798__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ net1440 net236 net397 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XANTENNA__10653__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ net881 top.a1.row1\[101\] _05114_ net891 vssd1 vssd1 vccd1 vccd1 _05166_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08631__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13030_ clknet_leaf_24_clk _00594_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10242_ net2070 net237 net454 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10173_ net243 net1987 net410 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
Xfanout1103 net1105 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_2
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input38_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout160 net163 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_2
Xfanout171 net174 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
XANTENNA__06970__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 _04764_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_1
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_199_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13863_ net1124 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__D_N _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06722__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12814_ clknet_leaf_115_clk _00378_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13794_ clknet_leaf_65_clk _01337_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08646__X _03757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12745_ clknet_leaf_3_clk _00309_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10828__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12676_ clknet_leaf_39_clk _00240_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06607__A _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _05460_ _05495_ _05452_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09424__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ _05368_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08822__A _01865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06789__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold608 top.DUT.register\[17\]\[31\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10509_ net158 net2282 net368 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__mux2_1
Xhold619 top.DUT.register\[16\]\[2\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10563__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ _05300_ _05333_ _05294_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a21o_1
XANTENNA__10990__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ clknet_leaf_9_clk _00792_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13159_ clknet_leaf_27_clk _00723_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09653__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06961__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ top.DUT.register\[9\]\[1\] net628 _02837_ _02844_ _02846_ vssd1 vssd1 vccd1
+ vccd1 _02847_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09372__B _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _02768_ _02769_ _02775_ _02777_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__or4_1
XANTENNA__09799__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ top.DUT.register\[9\]\[29\] net628 net605 top.DUT.register\[18\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
X_07582_ _02695_ _02705_ _02706_ _02708_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__or4_4
XFILLER_0_94_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13893__1143 vssd1 vssd1 vccd1 vccd1 _13893__1143/HI net1143 sky130_fd_sc_hd__conb_1
X_09321_ net907 top.pc\[15\] _04369_ net896 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__o211a_1
X_06533_ _01631_ _01634_ _01643_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__and3_1
XANTENNA__10738__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11423__A top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _02142_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06464_ top.a1.instruction\[22\] top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01591_ sky130_fd_sc_hd__and2_2
XFILLER_0_7_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07674__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ net313 _03297_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ net908 top.pc\[6\] _04240_ net898 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__o211a_1
X_06395_ _01496_ _01497_ net793 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__and3_2
XFILLER_0_172_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07426__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08134_ _03167_ _03176_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__or3b_2
XFILLER_0_71_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08065_ _01840_ net294 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__nand2_1
XANTENNA__10473__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_73_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout594_A _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ net1336 net865 _03031_ net593 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_A _01510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _03037_ _03039_ _03043_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__or4_2
XANTENNA__08179__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ net886 top.pc\[29\] net537 _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__a22o_1
XANTENNA__09850__X _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07849_ top.DUT.register\[16\]\[18\] net638 net622 top.DUT.register\[26\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06704__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10860_ net2189 net175 net349 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ top.a1.instruction\[27\] net822 _04540_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10791_ net2337 net193 net448 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
XANTENNA__10648__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ clknet_leaf_89_clk _00094_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07665__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12461_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[13\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[13\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_10_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11412_ _05246_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__or2_1
XANTENNA__07417__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ clknet_leaf_83_clk _00028_ net1014 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11343_ _05192_ _05194_ _01392_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__o21a_1
XANTENNA__10383__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06433__Y _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11274_ top.a1.row2\[27\] _05113_ _05117_ top.a1.row2\[11\] vssd1 vssd1 vccd1 vccd1
+ _05151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13013_ clknet_leaf_6_clk _00577_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ net171 net2310 net406 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__mux2_1
XANTENNA__07196__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net178 top.DUT.register\[8\]\[23\] net413 vssd1 vssd1 vccd1 vccd1 _00369_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06943__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09192__B _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ net185 net1992 net420 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XANTENNA__09893__A1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload3_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13846_ net1147 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_71_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13777_ clknet_leaf_64_clk _01320_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10558__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08448__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10989_ top.a1.data\[1\] top.a1.dataInTemp\[5\] net797 vssd1 vssd1 vccd1 vccd1 _05008_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12728_ clknet_leaf_109_clk _00292_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07120__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12659_ clknet_leaf_1_clk _00223_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06180_ top.a1.state\[2\] top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07439__Y _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 top.DUT.register\[31\]\[9\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10293__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold416 top.DUT.register\[22\]\[14\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__A2 _03715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 top.DUT.register\[12\]\[4\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 top.DUT.register\[23\]\[20\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold449 top.DUT.register\[6\]\[18\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout907 top.i_ready vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _04863_ _04864_ _04865_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a211o_1
Xfanout918 _01400_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07187__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout929 net933 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _01865_ _03921_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nand2_1
Xhold1105 top.DUT.register\[22\]\[24\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 top.DUT.register\[15\]\[25\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _03822_ _03856_ net277 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__mux2_1
Xhold1127 top.DUT.register\[20\]\[19\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 top.lcd.currentState\[3\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 top.DUT.register\[4\]\[9\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ _02820_ _02823_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nor3_4
XANTENNA__08136__B2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08683_ _02993_ _03338_ _03389_ _03770_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a221o_2
XANTENNA_fanout175_A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07634_ top.DUT.register\[20\]\[2\] net747 net674 top.DUT.register\[18\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07895__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07631__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10468__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ top.DUT.register\[3\]\[3\] net785 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__and2_1
XANTENNA__08439__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13849__1114 vssd1 vssd1 vccd1 vccd1 _13849__1114/HI net1114 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_192_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09304_ _01588_ _04352_ _04353_ net134 _04348_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout1084_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06516_ top.a1.instruction\[22\] top.a1.instruction\[23\] net801 vssd1 vssd1 vccd1
+ vccd1 _01643_ sky130_fd_sc_hd__and3b_2
XFILLER_0_152_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07647__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07496_ top.DUT.register\[20\]\[5\] net576 net556 top.DUT.register\[6\]\[5\] _02622_
+ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07111__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ _04270_ _04272_ _04271_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a21o_1
X_06447_ top.a1.instruction\[24\] top.a1.instruction\[27\] _01572_ _01573_ vssd1 vssd1
+ vccd1 vccd1 _01574_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout607_A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09166_ net133 _04217_ _04223_ _04224_ net908 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06378_ top.a1.instruction\[15\] top.a1.instruction\[16\] net810 vssd1 vssd1 vccd1
+ vccd1 _01505_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_32_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08117_ _03242_ _03243_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nand2_1
XANTENNA__10954__A0 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ _02739_ _02780_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09992__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ _03156_ _03160_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or2_2
Xhold950 top.DUT.register\[20\]\[28\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 top.DUT.register\[5\]\[29\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 top.DUT.register\[31\]\[8\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__C1 _03183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold983 top.DUT.register\[10\]\[20\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10931__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10706__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold994 top.DUT.register\[26\]\[3\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07178__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ net201 net1758 net427 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
XANTENNA__07365__X _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ net260 net1568 net425 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06925__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ _05796_ _05829_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_169_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ net231 net1565 net442 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XANTENNA__06689__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13700_ clknet_leaf_72_clk _01248_ net1096 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07886__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _05704_ _05737_ _05755_ _05761_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__a22oi_1
XANTENNA__07350__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ clknet_leaf_98_clk net1361 net982 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
X_10843_ net1810 net245 net352 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07638__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13562_ clknet_leaf_73_clk _01121_ net1093 vssd1 vssd1 vccd1 vccd1 top.a1.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ net1449 net257 net445 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08835__C1 _03935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06157__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ clknet_leaf_61_clk _00080_ net1099 vssd1 vssd1 vccd1 vccd1 top.ramstore\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_181_Right_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13493_ clknet_leaf_5_clk _01057_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11213__D net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12526__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12444_ clknet_leaf_95_clk top.ru.next_FetchedData\[28\] net991 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_152_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12375_ net2311 net117 _00017_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
XANTENNA__09187__B _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11326_ top.a1.dataIn\[26\] _05194_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__nor3_1
XANTENNA__07810__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892__1142 vssd1 vssd1 vccd1 vccd1 _13892__1142/HI net1142 sky130_fd_sc_hd__conb_1
XANTENNA__10841__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ top.a1.row2\[25\] _05113_ _05117_ top.a1.row2\[9\] _01444_ vssd1 vssd1 vccd1
+ vccd1 _05136_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07169__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10208_ net239 net2167 net405 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__mux2_1
X_11188_ net1224 net530 _05081_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__a21o_1
XANTENNA__06916__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ net243 net2020 net415 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07877__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13829_ clknet_leaf_68_clk _01370_ net1104 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10288__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ top.DUT.register\[13\]\[8\] net647 net564 top.DUT.register\[4\]\[8\] _02476_
+ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a221o_1
XANTENNA__07629__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08834__X _03935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06301_ top.lcd.currentState\[4\] _01445_ _01446_ top.lcd.nextState\[4\] vssd1 vssd1
+ vccd1 vccd1 _01448_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_174_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07281_ top.DUT.register\[28\]\[9\] net585 net690 top.DUT.register\[3\]\[9\] _02407_
+ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a221o_1
X_09020_ _03480_ _03508_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06232_ net1829 net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[8\] sky130_fd_sc_hd__and2_1
XANTENNA__09378__A top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08054__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06163_ top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XANTENNA__09097__B _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 top.ramload\[30\] vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09251__C1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold213 top.DUT.register\[19\]\[1\] vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09665__X _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 top.DUT.register\[23\]\[24\] vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold235 top.DUT.register\[7\]\[31\] vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 top.DUT.register\[29\]\[1\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 top.DUT.register\[16\]\[9\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 top.DUT.register\[13\]\[12\] vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 top.DUT.register\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ top.a1.instruction\[31\] _01622_ net527 _04913_ vssd1 vssd1 vccd1 vccd1 _04914_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10751__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 _01533_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 _01531_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_4
Xfanout726 _01525_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_8
X_09853_ _03915_ net343 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nand2_1
Xfanout737 _01521_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_8
Xfanout748 _01517_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 _01510_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06907__A2 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08804_ _03766_ _03905_ net312 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__mux2_1
XANTENNA__13055__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _04787_ _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__nand2_1
X_06996_ _01995_ _02037_ _02080_ _02121_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07580__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ _03765_ _03840_ net309 vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07632__Y _02759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09560__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _03774_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__nand2_2
XANTENNA__06529__X _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07332__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07617_ top.DUT.register\[11\]\[2\] net639 net556 top.DUT.register\[6\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
XANTENNA__10198__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ _02403_ _03708_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout724_A _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09987__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ top.DUT.register\[24\]\[4\] net737 net723 top.DUT.register\[14\]\[4\] _02664_
+ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10926__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ top.DUT.register\[28\]\[5\] net584 net674 top.DUT.register\[18\]\[5\] _02605_
+ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09218_ _04271_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ net233 net1464 net366 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12845__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09149_ net137 _04199_ _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07399__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ _06022_ _06026_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_112_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ net46 net857 vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10661__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__B _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ _05959_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__and2_1
Xhold780 top.DUT.register\[9\]\[4\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold791 top.DUT.register\[26\]\[5\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net22 net842 net812 net1324 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__o22a_1
XANTENNA__10233__Y _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07571__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12993_ clknet_leaf_25_clk _00557_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11944_ _05809_ _05810_ _05778_ _05803_ _05806_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_99_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11875_ _05699_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_123_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08086__B _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13614_ clknet_leaf_62_clk net1196 net1101 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
X_10826_ top.DUT.register\[28\]\[22\] net185 net356 vssd1 vssd1 vccd1 vccd1 _01008_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10757_ net213 net2098 net376 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13545_ clknet_leaf_4_clk _01109_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12082__A_N top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13476_ clknet_leaf_40_clk _01040_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10688_ net202 net1486 net379 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12427_ clknet_leaf_97_clk top.ru.next_FetchedData\[11\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12358_ top.pad.button_control.r_counter\[12\] top.pad.button_control.r_counter\[11\]
+ _06141_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__and3_1
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11309_ net1174 _01445_ _01446_ _05180_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10571__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] top.lcd.cnt_500hz\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__a31o_1
X_13848__1113 vssd1 vssd1 vccd1 vccd1 _13848__1113/HI net1113 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_52_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06350__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06850_ top.DUT.register\[20\]\[23\] net747 net696 top.DUT.register\[23\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XANTENNA__09661__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06781_ net516 _01905_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__nor2_1
XANTENNA__09839__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06770__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _02163_ net488 net520 _03632_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__o22a_1
XANTENNA__07314__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11110__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08451_ net472 _03554_ _03557_ net476 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__o22a_1
XFILLER_0_187_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07402_ top.DUT.register\[28\]\[7\] net652 net560 top.DUT.register\[23\]\[7\] _02528_
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a221o_1
XFILLER_0_175_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08382_ net319 _03498_ _03502_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07333_ _02453_ _02454_ _02455_ _02459_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10746__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout138_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ top.DUT.register\[31\]\[14\] net784 net780 top.DUT.register\[15\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09003_ _03526_ _04064_ _03554_ _03493_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__or4bb_1
X_06215_ wb.curr_state\[1\] wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__nor2_4
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07195_ top.DUT.register\[16\]\[15\] _01514_ net735 top.DUT.register\[24\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1047_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06589__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10481__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_clk_X clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _04896_ _04898_ net338 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_6_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout534 _01613_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_A _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _01665_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_4
Xfanout556 _01653_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_8
Xfanout567 _01649_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_4
X_09836_ _04834_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout578 _01633_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_8
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07553__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ top.DUT.register\[23\]\[20\] net562 net598 top.DUT.register\[27\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net802 _04773_ _04767_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__a21o_1
XANTENNA__06761__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ _03748_ _03824_ net304 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ net344 _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__or2_1
XANTENNA__08187__A _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_202_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07305__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08649_ _03075_ _03737_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_25_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11660_ _05487_ _05526_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__xnor2_1
X_13891__1141 vssd1 vssd1 vccd1 vccd1 _13891__1141/HI net1141 sky130_fd_sc_hd__conb_1
XFILLER_0_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10611_ net150 net2015 net389 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__mux2_1
XANTENNA__07069__A1 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _05452_ _05458_ _05459_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_115_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10656__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08634__B _03127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire913 _01408_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ clknet_leaf_51_clk _00894_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10542_ net1518 net156 net364 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__mux2_1
XANTENNA__06435__A _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13261_ clknet_leaf_23_clk _00825_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ net170 net1999 net370 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08569__A1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12212_ top.a1.row2\[43\] net845 net813 _05638_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__a22o_1
X_13192_ clknet_leaf_34_clk _00756_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ top.a1.dataIn\[2\] _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__and2b_1
XANTENNA__10391__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _05942_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__or2_1
X_11025_ net4 net841 net811 net1252 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__o22a_1
XANTENNA__08741__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06752__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08368__Y _03490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08097__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ clknet_leaf_121_clk _00540_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11235__B top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11927_ _05772_ _05791_ _05795_ _05771_ _05773_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11858_ _05722_ _05723_ _05725_ _05726_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10809_ net2092 net249 net353 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_106_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_103_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10566__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _05626_ _05629_ _05632_ _05638_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__or4bb_2
XTAP_TAPCELL_ROW_103_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ clknet_leaf_110_clk _01092_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07961__A_N net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08009__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__Y _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ clknet_leaf_1_clk _01023_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09757__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07783__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08980__B2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _02951_ _02993_ _03035_ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__or4b_1
XANTENNA__06991__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06902_ _02020_ _02022_ _02024_ _02028_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__or4_2
X_07882_ top.DUT.register\[11\]\[17\] net755 net681 top.DUT.register\[7\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09391__A top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__A2 _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09621_ _04643_ _04644_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__o21ai_1
X_06833_ top.DUT.register\[23\]\[23\] net560 net595 top.DUT.register\[27\]\[23\] _01959_
+ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a221o_1
XANTENNA__08732__B2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06743__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__B _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__A top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ net528 _04586_ _04423_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__o21a_2
X_06764_ top.DUT.register\[13\]\[25\] net648 net628 top.DUT.register\[9\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XANTENNA__12690__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ _02165_ _03618_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_65_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09483_ _01930_ _04508_ _04512_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06695_ top.DUT.register\[4\]\[26\] net768 net710 top.DUT.register\[9\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a22o_1
XFILLER_0_203_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ net1294 net838 net816 _03553_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ _02683_ _03450_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__nand2_1
XANTENNA__10476__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_A _04925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ top.DUT.register\[24\]\[9\] net549 net612 top.DUT.register\[14\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ _02732_ _02733_ _03418_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07247_ top.DUT.register\[27\]\[14\] net777 net734 top.DUT.register\[19\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09748__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06542__X _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ top.DUT.register\[23\]\[13\] net563 net605 top.DUT.register\[18\]\[13\] _02304_
+ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout889_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_2
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06982__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout342 _04684_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_4
Xfanout353 _04962_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_204_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout364 _04960_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 _04952_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_6
XANTENNA__07526__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _04945_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
X_09819_ net190 net1780 net439 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__mux2_1
Xfanout397 net400 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_8
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ clknet_leaf_14_clk _00394_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12761_ clknet_leaf_36_clk _00325_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ top.a1.dataIn\[2\] top.a1.dataIn\[3\] top.a1.dataIn\[0\] top.a1.dataIn\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_120_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ clknet_leaf_45_clk _00256_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13847__1112 vssd1 vssd1 vccd1 vccd1 _13847__1112/HI net1112 sky130_fd_sc_hd__conb_1
X_11643_ _05465_ _05491_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__xor2_2
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10386__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _05441_ _05442_ top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06165__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_10525_ net1846 net219 net364 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__mux2_1
Xinput39 nrst vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_4
X_13313_ clknet_leaf_27_clk _00877_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09739__A0 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09476__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ clknet_leaf_55_clk _00808_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ net235 net2051 net369 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XANTENNA__08380__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ clknet_leaf_77_clk _00739_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10387_ net246 net1988 net327 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
X_12126_ _05983_ _05995_ _05979_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a21o_1
XANTENNA__07765__A2 _02543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__B2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06973__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _05905_ _05922_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11008_ top.a1.dataIn\[11\] net848 net843 _05020_ vssd1 vssd1 vccd1 vccd1 _05021_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output51_A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09911__B1 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__B2 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06725__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12959_ clknet_leaf_115_clk _00523_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06480_ _01580_ net902 net820 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__or3b_2
XFILLER_0_87_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10296__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08150_ net292 _02970_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11218__A_N net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07101_ top.DUT.register\[28\]\[10\] net651 net595 top.DUT.register\[27\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08081_ _02099_ net295 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07032_ top.DUT.register\[28\]\[11\] net653 net622 top.DUT.register\[26\]\[11\] _02148_
+ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a221o_1
XANTENNA__07458__X _02585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08290__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__A _01929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_184_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ top.pc\[1\] _02788_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nand2_1
XANTENNA__06964__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890__1140 vssd1 vssd1 vccd1 vccd1 _13890__1140/HI net1140 sky130_fd_sc_hd__conb_1
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ top.DUT.register\[11\]\[16\] net640 net620 top.DUT.register\[26\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_149_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08289__X _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07865_ _02970_ _02990_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__and2_1
XANTENNA__06716__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_A _04958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12463__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _04629_ net847 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__nor2_1
X_06816_ _01936_ _01937_ _01939_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_162_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ top.DUT.register\[28\]\[19\] net586 net741 top.DUT.register\[8\]\[19\] _02922_
+ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a221o_1
XANTENNA__06192__B2 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09535_ top.pc\[28\] _04557_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or2_1
X_06747_ _01867_ _01868_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__or3_1
XANTENNA__08469__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_A _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ top.pc\[24\] _04483_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_195_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06537__X _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06678_ top.DUT.register\[9\]\[27\] net627 _01802_ _01803_ _01804_ vssd1 vssd1 vccd1
+ vccd1 _01805_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_195_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07141__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ _03425_ _03536_ net308 vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__mux2_2
XFILLER_0_191_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ _04439_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08348_ _03467_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12143__A_N top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08279_ _03267_ _03286_ net286 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux2_1
XANTENNA__10934__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ net1437 net239 net397 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XANTENNA__07995__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net1216 net824 _05165_ net1095 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ net1774 net239 net454 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10172_ net248 net1688 net409 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
XANTENNA__06955__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_4
Xfanout150 _04691_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout161 net163 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
Xfanout172 net173 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_2
Xfanout183 net186 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_2
Xfanout194 _04811_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06707__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13862_ net1123 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08927__X _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11059__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ clknet_leaf_23_clk _00377_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13793_ clknet_leaf_65_clk _01336_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12744_ clknet_leaf_35_clk _00308_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_177_Left_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07132__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07683__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ clknet_leaf_33_clk _00239_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ _05460_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ _05388_ _05395_ _05397_ net250 _05392_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a41o_1
XANTENNA__10844__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08632__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07986__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold609 top.DUT.register\[25\]\[28\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ net161 net1892 net365 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__mux2_1
X_11488_ _05294_ _05300_ net267 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__nand3_1
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10990__A1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10439_ net173 net1296 net325 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__mux2_1
X_13227_ clknet_leaf_29_clk _00791_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_186_Left_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07199__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08935__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ clknet_leaf_24_clk _00722_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06946__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ _05966_ _05967_ _05975_ _05972_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a31o_1
X_13089_ clknet_leaf_25_clk _00653_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11298__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07650_ top.DUT.register\[26\]\[2\] net759 net704 top.DUT.register\[15\]\[2\] _02776_
+ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_195_Right_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07371__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06601_ top.DUT.register\[4\]\[29\] net565 net601 top.DUT.register\[10\]\[29\] _01727_
+ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a221o_1
XANTENNA__07910__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ top.DUT.register\[2\]\[3\] net659 net552 top.DUT.register\[7\]\[3\] _02707_
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ net136 _04356_ _04368_ net907 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07460__Y _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06532_ net900 _01592_ net801 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__and3_2
XANTENNA__08285__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07123__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ _01615_ _02210_ _04303_ net823 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_177_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06463_ top.a1.instruction\[20\] top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ _01590_ sky130_fd_sc_hd__and2_2
XFILLER_0_173_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08871__B1 _03963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08202_ net316 _03327_ _03312_ net272 vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__X _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ net137 _04227_ _04239_ net908 vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__o211ai_1
X_06394_ _01498_ net792 _01505_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__and3_4
X_08133_ net481 _03190_ _03254_ _03259_ _03181_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08623__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10754__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout218_A _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10430__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_08064_ _01797_ net291 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _02131_ _02136_ _02141_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__or3_4
XFILLER_0_12_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_4__f_clk_X clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06937__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06401__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ net1256 net870 _03072_ net593 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__a22o_1
X_07917_ top.DUT.register\[23\]\[16\] net696 net675 top.DUT.register\[18\]\[16\] _03040_
+ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08897_ _03974_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout754_A _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_197_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ top.DUT.register\[17\]\[18\] net646 net559 top.DUT.register\[6\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__a22o_1
XANTENNA__11317__C top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07362__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07901__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10929__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _02905_ _02165_ _02162_ _02143_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08466__Y _03584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ top.pc\[27\] _04532_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__xnor2_1
X_10790_ net1747 net204 net447 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__mux2_1
XANTENNA__08195__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08963__A1_N net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ _04472_ _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ clknet_leaf_96_clk top.ru.next_FetchedInstr\[12\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ _05245_ _05275_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10664__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ clknet_leaf_83_clk _00027_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08978__A1_N net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ _05203_ _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06640__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ top.a1.row1\[107\] _05116_ _05118_ top.a1.row2\[19\] _05149_ vssd1 vssd1
+ vccd1 vccd1 _05150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13012_ clknet_leaf_59_clk _00576_ net1109 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10224_ net177 net2273 net405 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10155_ net186 net1559 net415 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10086_ net188 net2039 net419 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
Xhold6 top.ramaddr\[23\] vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08089__B _03012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07353__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13845_ net1146 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10839__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_15__f_clk_X clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__A0 _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13776_ clknet_leaf_65_clk _01319_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10988_ net1455 _05007_ net535 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
XANTENNA__08448__A3 _03565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12727_ clknet_leaf_105_clk _00291_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ clknet_leaf_51_clk _00222_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _05475_ _05477_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10574__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12589_ clknet_leaf_32_clk _00153_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_194_Left_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold406 top.DUT.register\[9\]\[18\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10963__A1 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 top.DUT.register\[23\]\[27\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap125 _06029_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
Xhold428 top.DUT.register\[5\]\[9\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 top.DUT.register\[28\]\[8\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13257__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06631__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06919__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net910 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_2
Xfanout919 net934 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03885_ _03920_ _01907_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_14__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__07592__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 top.DUT.register\[13\]\[28\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 top.DUT.register\[20\]\[15\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _03205_ _03209_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__nand2_1
Xhold1128 top.DUT.register\[19\]\[10\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1139 top.DUT.register\[10\]\[17\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__C1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07702_ _02824_ _02826_ _02828_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__or3_2
XFILLER_0_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08682_ _02992_ net488 net486 _02991_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_wire510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06698__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ net806 _02739_ _02758_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__o21a_1
XANTENNA__10749__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout168_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ _02690_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__inv_2
XANTENNA__07631__B _02757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_192_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06515_ _01591_ _01631_ _01634_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__and3_4
X_09303_ _04350_ _04351_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07495_ top.DUT.register\[30\]\[5\] net615 net544 top.DUT.register\[5\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06446_ top.a1.instruction\[22\] top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01573_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _04286_ _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ _04218_ _04222_ _01619_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__a21o_1
XANTENNA__06870__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06377_ top.a1.instruction\[19\] _01498_ _01503_ vssd1 vssd1 vccd1 vccd1 _01504_
+ sky130_fd_sc_hd__and3_4
XANTENNA__10484__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06534__Y _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ _02298_ net290 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09096_ _04156_ _04157_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08047_ _03164_ _03172_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__or2_1
Xhold940 top.DUT.register\[22\]\[11\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold951 top.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 top.DUT.register\[21\]\[16\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 top.DUT.register\[20\]\[16\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 top.DUT.register\[15\]\[21\] vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 top.DUT.register\[4\]\[19\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ net266 top.DUT.register\[4\]\[1\] net426 vssd1 vssd1 vccd1 vccd1 _00219_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_209_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ net34 top.ru.state\[0\] _01429_ _01484_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_68_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _05822_ _05823_ _05796_ _05801_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a211o_1
XANTENNA__07335__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07822__A _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ net238 net2132 net441 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07886__A1 top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06689__A2 _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _05656_ _05701_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__xnor2_1
X_13630_ clknet_leaf_61_clk net1223 net1100 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
X_10842_ net1412 net246 net349 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13561_ clknet_leaf_69_clk top.a1.nextHex\[4\] net1103 vssd1 vssd1 vccd1 vccd1 _01381_
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10773_ net1488 net260 net445 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12512_ clknet_leaf_61_clk _00079_ net1101 vssd1 vssd1 vccd1 vccd1 top.ramstore\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13492_ clknet_leaf_61_clk _01056_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ clknet_leaf_95_clk top.ru.next_FetchedData\[27\] net990 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[27\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__10394__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06861__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12374_ net2202 net912 net38 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06613__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ _05185_ _05192_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11256_ top.a1.row1\[121\] _05106_ _05116_ top.a1.row1\[105\] _05134_ vssd1 vssd1
+ vccd1 vccd1 _05135_ sky130_fd_sc_hd__a221o_1
XANTENNA__08543__B1_N _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ net244 net2109 net408 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__mux2_1
X_11187_ net850 _05067_ net531 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07574__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ net249 net1863 net413 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_59_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_128_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ net253 net1695 net419 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11122__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07326__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10569__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13828_ clknet_leaf_69_clk net1173 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13759_ clknet_leaf_74_clk _01302_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_06300_ _01447_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07280_ top.DUT.register\[18\]\[9\] net675 _02405_ _02406_ vssd1 vssd1 vccd1 vccd1
+ _02407_ sky130_fd_sc_hd__a211o_1
XANTENNA__06301__B2 top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06231_ net1415 net873 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[7\] sky130_fd_sc_hd__and2_1
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06852__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06162_ top.a1.dataIn\[24\] vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold203 top.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 top.a1.data\[5\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 top.DUT.register\[28\]\[9\] vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 top.DUT.register\[27\]\[1\] vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold247 top.DUT.register\[27\]\[14\] vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 top.DUT.register\[7\]\[9\] vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 top.DUT.register\[29\]\[20\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net835 _04623_ _04911_ _01586_ _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o221ai_1
XANTENNA__07907__A _03012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 _01533_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_2
XFILLER_0_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout716 net719 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_8
Xfanout727 _01523_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_8
X_09852_ net173 net1561 net439 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__mux2_1
Xfanout738 _01521_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
Xfanout749 _01517_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_8
X_08803_ _03840_ _03904_ net307 vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__mux2_1
X_09783_ top.pc\[18\] _04407_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__or2_1
X_06995_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout285_A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09306__A1 top.i_ready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _03800_ _03839_ net282 vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07317__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _03033_ net489 net474 _03760_ _03769_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o221a_1
XANTENNA__10479__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ top.DUT.register\[29\]\[2\] net663 net611 top.DUT.register\[14\]\[2\] _02742_
+ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a221o_1
X_08596_ _02403_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_159_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07547_ _02666_ _02668_ _02670_ _02673_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__or4_1
XANTENNA__08817__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout717_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07478_ top.DUT.register\[4\]\[5\] net767 net704 top.DUT.register\[15\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XANTENNA__07096__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09217_ _02423_ _02427_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__or2_1
XANTENNA__06843__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06429_ top.DUT.register\[21\]\[30\] net693 net671 top.DUT.register\[16\]\[30\] _01555_
+ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09148_ net133 _04204_ _04206_ _04207_ net910 vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09079_ _04137_ _04138_ _04139_ _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_112_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11110_ net917 net1555 net852 _05041_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a31o_1
XFILLER_0_188_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ _05935_ _05937_ _05945_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__mux2_1
Xhold770 top.DUT.register\[24\]\[12\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 top.DUT.register\[31\]\[26\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold792 top.DUT.register\[17\]\[18\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11041_ net21 net842 net812 net1325 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__o22a_1
XANTENNA__06440__B net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ clknet_leaf_47_clk _00556_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11943_ _05805_ _05807_ _05811_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__and3b_1
XANTENNA__10389__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08520__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06168__A top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11874_ _05695_ _05704_ net131 _05701_ _05656_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_123_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ clknet_leaf_114_clk net1236 net939 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10825_ net1405 net189 net356 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13544_ clknet_leaf_35_clk _01108_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07087__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10756_ net217 net1842 net373 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13475_ clknet_leaf_50_clk _01039_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06834__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ net210 net1930 net378 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
X_12426_ clknet_leaf_97_clk top.ru.next_FetchedData\[10\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12357_ _06142_ _06143_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10852__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ _05093_ _05096_ _05103_ _05177_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a211oi_1
X_12288_ _01437_ _06098_ _06100_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__and3_1
X_11239_ net884 _05093_ net882 vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_52_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07011__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13535__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06780_ net516 _01905_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07462__A _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10299__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08450_ net479 _03560_ _03566_ net519 _03568_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__o221a_1
X_07401_ top.DUT.register\[6\]\[7\] net556 net611 top.DUT.register\[14\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a22o_1
X_08381_ net270 _03499_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07332_ top.DUT.register\[15\]\[8\] net704 net689 top.DUT.register\[3\]\[8\] _02457_
+ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a221o_1
XANTENNA__11712__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12488__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ top.DUT.register\[8\]\[14\] net569 net602 top.DUT.register\[10\]\[14\] _02389_
+ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09002_ _03416_ _03449_ _04063_ _03465_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__or4b_1
X_06214_ net34 net865 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08580__X _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ top.DUT.register\[22\]\[15\] net752 net681 top.DUT.register\[7\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a22o_1
XANTENNA__10762__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout200_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07786__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ net804 _04894_ _04895_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a31o_1
Xfanout524 _01617_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07538__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout535 _04989_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07002__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ top.pc\[23\] _04493_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__or2_1
Xfanout557 _01653_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
Xfanout568 net571 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_8
Xfanout579 _01633_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _04768_ _04771_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__xnor2_1
X_06978_ top.DUT.register\[29\]\[20\] net666 net546 top.DUT.register\[5\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a22o_1
X_08717_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout834_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ top.a1.dataIn\[7\] net794 net803 top.pc\[7\] _04712_ vssd1 vssd1 vccd1 vccd1
+ _04713_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_202_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ net1273 net839 net818 _03758_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a22o_1
XANTENNA__08755__X _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _02403_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10610_ net142 net1853 net387 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08266__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _05458_ _05459_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net2056 net161 net361 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06435__B _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13260_ clknet_leaf_10_clk _00824_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ net171 net1845 net370 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
X_12211_ top.a1.row2\[42\] net845 net813 _05677_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__a22o_1
XANTENNA__10672__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ clknet_leaf_7_clk _00755_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ _05992_ _06001_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07241__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12073_ _05912_ _05923_ _05927_ _05925_ _05924_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__a311o_1
XANTENNA__07529__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ net3 net831 net830 net2111 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__a22o_1
XANTENNA__09481__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12975_ clknet_leaf_51_clk _00539_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11926_ _05772_ _05791_ _05795_ _05771_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a22o_2
XFILLER_0_185_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07701__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11857_ _05725_ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__nand2_2
XANTENNA__10847__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ net2319 net251 net355 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__mux2_1
XANTENNA__08257__A1 _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08257__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ _05653_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13527_ clknet_leaf_16_clk _01091_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06807__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ net150 net1667 net373 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13458_ clknet_leaf_48_clk _01022_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12409_ clknet_leaf_88_clk _00045_ net1005 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10582__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
X_13389_ clknet_leaf_23_clk _00953_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07950_ _03075_ _03076_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__or2_2
XANTENNA__06991__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ top.DUT.register\[1\]\[22\] net658 _02018_ _02025_ _02027_ vssd1 vssd1 vccd1
+ vccd1 _02028_ sky130_fd_sc_hd__a2111o_1
X_07881_ top.DUT.register\[19\]\[17\] net731 net685 top.DUT.register\[1\]\[17\] _03007_
+ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_182_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08559__Y _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _04645_ _04646_ _04647_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__o22a_1
XANTENNA__08732__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ top.DUT.register\[29\]\[23\] net663 net607 top.DUT.register\[12\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a22o_1
XANTENNA__07940__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__A _02298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ top.a1.instruction\[29\] net821 _04540_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__o21a_1
X_06763_ top.DUT.register\[5\]\[25\] net545 net596 top.DUT.register\[27\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
X_08502_ _02235_ _03595_ _02905_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09482_ _04519_ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06694_ _01818_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_65_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12669__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08433_ net887 top.pc\[7\] net538 _03552_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10757__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout150_A _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08248__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08364_ net519 _03475_ _03485_ net479 _03482_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07315_ top.DUT.register\[21\]\[9\] net572 net600 top.DUT.register\[10\]\[9\] _02441_
+ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08295_ _03415_ _03418_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07246_ top.DUT.register\[12\]\[14\] net582 net698 top.DUT.register\[23\]\[14\] _02372_
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a221o_1
XANTENNA__07471__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09748__A1 _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07177_ top.DUT.register\[26\]\[13\] net621 net597 top.DUT.register\[27\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07367__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08420__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__Y _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout784_A _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06431__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout310 net312 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_167_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_4
Xfanout332 net333 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
Xfanout343 _04683_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_4
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 _04962_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_204_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout365 _04959_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_6
Xfanout376 _04952_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
X_09818_ _03847_ net340 net337 _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__o211a_4
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
Xfanout398 net400 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_6
XANTENNA__08198__A _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09749_ net195 net1460 net439 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12760_ clknet_leaf_13_clk _00324_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09684__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11711_ _05530_ _05559_ _05573_ _05580_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_120_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ clknet_leaf_1_clk _00255_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10667__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11642_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08239__B2 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06446__A top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11573_ _05441_ _05442_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08932__Y _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ clknet_leaf_44_clk _00876_ net1080 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ net2288 net223 net361 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ clknet_leaf_47_clk _00807_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09476__B top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ net241 net1908 net370 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08380__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ clknet_leaf_121_clk _00738_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07214__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10386_ net253 net2058 net329 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
X_12125_ _05967_ _05982_ _05975_ _05974_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_176_Right_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12056_ _05924_ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ top.a1.data\[7\] top.a1.dataInTemp\[11\] net797 vssd1 vssd1 vccd1 vccd1 _05020_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08714__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07922__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output44_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12958_ clknet_leaf_13_clk _00522_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09675__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11909_ _05740_ _05758_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_47_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10577__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ clknet_leaf_37_clk _00453_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__B1 top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07100_ top.DUT.register\[4\]\[10\] net567 net545 top.DUT.register\[5\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XANTENNA__07989__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ _03205_ _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07031_ _02151_ _02153_ _02154_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06661__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08290__B _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07205__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08402__B2 _03522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ _01386_ net896 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ top.DUT.register\[29\]\[16\] net664 net648 top.DUT.register\[13\]\[16\] _03059_
+ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout198_A _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _02970_ _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__nor2_1
XANTENNA__07913__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ top.a1.state\[1\] net893 top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04635_
+ sky130_fd_sc_hd__or3b_1
X_06815_ top.DUT.register\[23\]\[24\] net563 net605 top.DUT.register\[18\]\[24\] _01941_
+ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ top.DUT.register\[14\]\[19\] net723 net672 top.DUT.register\[16\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout365_A _04959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ top.pc\[28\] _04557_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06746_ top.DUT.register\[25\]\[25\] net771 net581 top.DUT.register\[12\]\[25\] _01872_
+ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10487__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _04501_ _04502_ _04503_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06677_ top.DUT.register\[16\]\[27\] net635 net548 top.DUT.register\[24\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_195_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12432__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08416_ _03476_ _03535_ net281 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07692__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ top.pc\[20\] _04425_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08347_ _03409_ _03468_ net311 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07444__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ net269 _03401_ _03398_ net270 vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_78_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout999_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06652__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07229_ top.DUT.register\[18\]\[15\] net603 net540 top.DUT.register\[22\]\[15\] _02355_
+ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a221o_1
XANTENNA__09296__B _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ net2326 net244 net456 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net251 net1940 net410 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout140 net143 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_2
Xfanout151 _04691_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_2
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_98_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout195 net198 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
X_13861_ net1122 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12812_ clknet_leaf_11_clk _00376_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13792_ clknet_leaf_67_clk _01335_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12743_ clknet_leaf_7_clk _00307_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10397__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12674_ clknet_leaf_43_clk _00238_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06176__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07683__A2 _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06891__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _05449_ _05461_ _05480_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_100_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11232__D net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11810__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09487__A top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11556_ _05388_ _05397_ net250 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06643__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10507_ net164 net2112 net368 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11487_ _05355_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10990__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_40_clk _00790_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10438_ net177 net1761 net323 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12414__Q top.i_ready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ clknet_leaf_119_clk _00721_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10860__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10369_ net466 _04926_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nand2_8
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12108_ _05966_ _05967_ _05975_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__and3_1
X_13088_ clknet_leaf_46_clk _00652_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12039_ _05886_ _05908_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06600_ top.DUT.register\[23\]\[29\] net562 net553 top.DUT.register\[7\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07580_ top.DUT.register\[25\]\[3\] net624 net607 top.DUT.register\[12\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire500_A _02469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06531_ top.DUT.register\[3\]\[30\] net786 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08285__B _03127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10100__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ net529 _02734_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__or2_1
X_06462_ net903 _01494_ _01584_ _01587_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08853__X _03953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08871__A1 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07674__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ net300 _03326_ _03319_ net285 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06882__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06393_ _01496_ net793 _01503_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__and3_4
X_09181_ net133 _04232_ _04238_ net819 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__o22a_1
X_08132_ _03256_ _03257_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__nor2_2
XFILLER_0_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07426__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09382__A_N _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06634__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07014_ _02126_ _02127_ _02139_ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__or4_1
XANTENNA__09684__X _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10194__A0 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10770__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1022_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ net504 net591 net1177 net867 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout482_A _03184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ top.DUT.register\[12\]\[16\] net581 net736 top.DUT.register\[24\]\[16\] _03042_
+ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a221o_1
X_08896_ _03990_ _03993_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__nor2_2
X_07847_ top.DUT.register\[25\]\[18\] net626 net613 top.DUT.register\[14\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_197_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__D top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A2_N _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07778_ _02184_ _02232_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__and2b_1
XFILLER_0_195_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _04552_ _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06729_ top.DUT.register\[6\]\[26\] net559 net618 top.DUT.register\[30\]\[26\] _01845_
+ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout914_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10010__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ _04471_ _04473_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__nand2_1
XANTENNA__07665__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06873__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ _01622_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ _05241_ _05266_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__xor2_2
XFILLER_0_105_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07417__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ clknet_leaf_88_clk _00026_ net1005 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06625__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _05205_ _05210_ _05209_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a21boi_1
XANTENNA__13401__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06443__B _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11272_ top.a1.row1\[3\] _05094_ _05111_ top.a1.row2\[3\] vssd1 vssd1 vccd1 vccd1
+ _05149_ sky130_fd_sc_hd__a22o_1
XANTENNA__13059__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ clknet_leaf_1_clk _00575_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10223_ net184 net1614 net408 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__mux2_1
XANTENNA__10680__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07050__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ net187 net1730 net415 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold7 top.lcd.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net193 top.DUT.register\[6\]\[20\] net420 vssd1 vssd1 vccd1 vccd1 _00302_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09878__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13844_ net1145 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13775_ clknet_leaf_65_clk _01318_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07105__A1 _02231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ top.a1.dataIn\[4\] net848 net843 _05006_ vssd1 vssd1 vccd1 vccd1 _05007_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12726_ clknet_leaf_120_clk _00290_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08853__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10855__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12657_ clknet_leaf_3_clk _00221_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12588_ clknet_leaf_11_clk _00152_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06616__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ _01393_ _05407_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__xnor2_2
Xhold407 top.DUT.register\[18\]\[12\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap126 _05988_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold429 top.DUT.register\[29\]\[10\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08369__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13209_ clknet_leaf_36_clk _00773_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10590__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_55_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07041__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08750_ _03507_ _03541_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__nand2_1
Xhold1107 top.DUT.register\[12\]\[8\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 top.DUT.register\[5\]\[27\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 top.DUT.register\[22\]\[23\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__X _02879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ top.DUT.register\[8\]\[0\] net739 net671 top.DUT.register\[16\]\[0\] _02827_
+ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a221o_1
X_08681_ net273 _03788_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07344__A1 top.a1.instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__B1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07632_ net806 _02739_ _02758_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_179_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ top.a1.instruction\[24\] net528 _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a21oi_2
X_09302_ _04350_ _04351_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__nor2_1
X_06514_ _01632_ _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__nor2_4
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09679__X _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07647__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ top.DUT.register\[21\]\[5\] net572 net552 top.DUT.register\[7\]\[5\] _02620_
+ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _02184_ _02212_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__nand2_1
XANTENNA__10765__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06445_ top.a1.instruction\[28\] top.a1.instruction\[29\] top.a1.instruction\[30\]
+ top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout328_A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09164_ _04218_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nor2_1
X_06376_ top.a1.instruction\[16\] net810 top.a1.instruction\[15\] vssd1 vssd1 vccd1
+ vccd1 _01503_ sky130_fd_sc_hd__and3b_2
XANTENNA__10939__C1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ net506 net295 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09095_ _02835_ net494 vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08046_ _03164_ _03172_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_170_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold930 top.pad.button_control.r_counter\[13\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 top.DUT.register\[22\]\[27\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold952 top.DUT.register\[18\]\[26\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 top.DUT.register\[25\]\[13\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 top.lcd.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 top.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 top.ramload\[20\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09997_ net150 net1859 net425 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ net865 _01483_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__or2_4
XANTENNA__10005__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ net1247 net839 net817 _03977_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ net239 net2219 net441 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ net129 _05749_ _05757_ _05740_ _05735_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07886__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10841_ net2343 net254 net351 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ clknet_leaf_69_clk top.a1.nextHex\[3\] net1103 vssd1 vssd1 vccd1 vccd1 _01380_
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07638__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08835__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ net1396 net264 net447 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08835__B2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ clknet_leaf_114_clk _00078_ net939 vssd1 vssd1 vccd1 vccd1 top.ramstore\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06846__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10675__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ clknet_leaf_1_clk _01055_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ clknet_leaf_95_clk top.ru.next_FetchedData\[26\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12373_ net2188 net912 net37 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11324_ _05189_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__and2_2
XANTENNA__07810__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11255_ top.a1.row1\[1\] _05094_ _05120_ top.a1.row2\[41\] vssd1 vssd1 vccd1 vccd1
+ _05134_ sky130_fd_sc_hd__a22o_1
XANTENNA__06460__Y _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ net248 net2023 net405 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11186_ net1204 net530 _05080_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__a21o_1
X_10137_ net251 net1318 net415 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ net255 net2240 net417 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__mux2_1
XANTENNA__08387__Y _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__B1 _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07877__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13827_ clknet_leaf_69_clk _01368_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_35_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07629__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ clknet_leaf_73_clk _01301_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12709_ clknet_leaf_117_clk _00273_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06837__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13689_ clknet_leaf_74_clk _01237_ net1088 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06301__A2 _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06230_ top.ramload\[6\] net874 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[6\]
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06161_ top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 top.DUT.register\[27\]\[21\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold215 top.DUT.register\[14\]\[16\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold226 top.ramload\[18\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold237 top.DUT.register\[11\]\[13\] vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ top.a1.dataIn\[31\] net332 net334 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a21oi_2
Xhold248 top.DUT.register\[29\]\[15\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold259 top.DUT.register\[6\]\[9\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout706 _01533_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_6
Xfanout717 net718 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ net336 _04841_ _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and3_2
Xfanout728 _01523_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
Xfanout739 _01519_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
X_08802_ _03872_ _03903_ net281 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__mux2_1
X_09782_ top.pc\[18\] _04407_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11148__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06994_ _02119_ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08733_ _03268_ _03273_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout180_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08664_ net472 _03762_ _03763_ net521 _03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__o221a_1
XANTENNA__07868__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07615_ top.DUT.register\[17\]\[2\] net643 net599 top.DUT.register\[10\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08595_ _03664_ _03707_ _02318_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout445_A _04950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ top.DUT.register\[8\]\[4\] net741 net724 top.DUT.register\[17\]\[4\] _02672_
+ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a221o_1
XANTENNA__08817__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06828__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ top.DUT.register\[30\]\[5\] net712 net681 top.DUT.register\[7\]\[5\] _02603_
+ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout612_A _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13810__D _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ _02423_ _02427_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__and2_1
X_06428_ top.DUT.register\[20\]\[30\] net748 net668 top.DUT.register\[5\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09147_ _04192_ _04195_ _04205_ _01619_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__a31o_1
X_06359_ net904 top.a1.instruction\[6\] _01475_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ _01694_ _01736_ _01953_ _03152_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08029_ _01569_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__nand2_1
Xhold760 top.DUT.register\[29\]\[24\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 top.DUT.register\[25\]\[2\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold782 top.DUT.register\[14\]\[21\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net20 net832 _05024_ net1675 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold793 top.DUT.register\[17\]\[22\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10560__A0 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12991_ clknet_leaf_115_clk _00555_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_71_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__inv_2
XANTENNA__06449__A top.a1.instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__Y _03127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13834__RESET_B net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11873_ _05707_ _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_28_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ clknet_leaf_75_clk net1275 net1090 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ net1918 net191 net355 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13543_ clknet_leaf_7_clk _01107_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06819__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11812__B1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ net227 net1839 net374 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13474_ clknet_leaf_44_clk _01038_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07492__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ net220 net2074 net380 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_80_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ clknet_leaf_97_clk top.ru.next_FetchedData\[9\] net984 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_180_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12356_ net1843 _06141_ net796 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06598__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ net1212 _01443_ _05179_ net1095 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__o211a_1
X_12287_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__a21o_1
X_11238_ net882 net884 _05109_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12422__Q top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ net1353 net532 net525 _05072_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06770__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06359__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ top.DUT.register\[30\]\[7\] net616 net544 top.DUT.register\[5\]\[7\] _02523_
+ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ net316 net285 _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12614__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07331_ top.DUT.register\[12\]\[8\] net580 net751 top.DUT.register\[22\]\[8\] _02456_
+ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a221o_1
XANTENNA__11712__B top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07262_ top.DUT.register\[13\]\[14\] net649 net614 top.DUT.register\[14\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09001_ _02881_ _03168_ net473 _02783_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__or4b_1
XFILLER_0_155_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06213_ net866 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07193_ _02318_ _02319_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__nor2_2
XFILLER_0_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07235__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06589__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ _04587_ net526 net332 top.a1.dataIn\[29\] net334 vssd1 vssd1 vccd1 vccd1
+ _04897_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout525 _05065_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout536 net538 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ top.pc\[23\] _04493_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__nand2_1
Xfanout547 _01665_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1102_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 _01653_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_8
Xfanout569 net571 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_206_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ _04771_ _04768_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__and2b_1
X_06977_ top.DUT.register\[12\]\[20\] net610 net606 top.DUT.register\[18\]\[20\] _02103_
+ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout562_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _03786_ _03822_ net277 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XANTENNA__11098__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09696_ net836 _04243_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__nor2_1
XANTENNA__09316__A_N _02339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08647_ net886 top.pc\[16\] net539 _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _02899_ _03669_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07529_ top.DUT.register\[29\]\[4\] net666 net654 top.DUT.register\[28\]\[4\] _02655_
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a221o_1
XFILLER_0_181_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ net1712 net165 net364 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__mux2_1
XANTENNA__11270__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07474__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08771__X _03875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10471_ net176 net1651 net369 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12210_ top.a1.row2\[41\] net845 net813 net130 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07226__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ clknet_leaf_19_clk _00754_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ _06004_ _06007_ _06008_ _06010_ _05999_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__o32a_2
XTAP_TAPCELL_ROW_94_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12072_ _05916_ _05930_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold590 top.DUT.register\[31\]\[0\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08726__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net33 net841 net811 net1302 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__o22a_1
XANTENNA__08659__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06752__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12974_ clknet_leaf_116_clk _00538_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_X clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ _05770_ _05787_ _05789_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__or3_2
XFILLER_0_197_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11813__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11856_ _05685_ net130 _05686_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a21o_1
XFILLER_0_196_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10807_ net1443 net255 net353 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_109_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11787_ _05632_ _05654_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__and3_1
XANTENNA__08257__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11261__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13526_ clknet_leaf_2_clk _01090_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07465__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10738_ net142 net1893 net383 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12417__Q top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ clknet_leaf_118_clk _01021_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09206__A1 _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ net1900 net164 net452 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07217__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ clknet_leaf_89_clk _00044_ net1006 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12210__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_8_clk _00952_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_12339_ top.pad.button_control.r_counter\[5\] top.pad.button_control.r_counter\[4\]
+ _06128_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06900_ top.DUT.register\[13\]\[22\] net649 net543 top.DUT.register\[22\]\[22\] _02026_
+ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a221o_1
XANTENNA__06991__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ top.DUT.register\[31\]\[17\] net743 net678 top.DUT.register\[13\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_182_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06831_ top.DUT.register\[2\]\[23\] net659 net655 top.DUT.register\[1\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a22o_1
XANTENNA__06743__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ top.pc\[29\] _04566_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10103__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ top.DUT.register\[12\]\[25\] net608 net603 top.DUT.register\[18\]\[25\] _01888_
+ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a221o_1
X_08501_ net1347 net838 net817 _03617_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09481_ _04518_ net517 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_65_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06693_ _01797_ _01816_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__nor2_1
XANTENNA__08575__Y _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08432_ _03334_ _03526_ _03551_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ net320 _03484_ _03474_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_92_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08248__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout143_A _04915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07314_ top.DUT.register\[2\]\[9\] net660 net620 top.DUT.register\[26\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a22o_1
XANTENNA__07456__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__A1 top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__X _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _02783_ _03379_ _02781_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_190_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ top.DUT.register\[29\]\[14\] net702 net683 top.DUT.register\[7\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout310_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10773__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1052_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07208__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09748__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ top.DUT.register\[1\]\[13\] net657 net558 top.DUT.register\[6\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
XANTENNA__08956__B1 _02585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07367__B _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06982__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11307__A2 _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 _02662_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_4
Xfanout333 _04766_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_2
Xfanout344 _04683_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
Xfanout355 _04962_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_6
Xfanout366 _04959_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
Xfanout377 _04949_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_6
X_09817_ net802 _04815_ _04816_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a31o_1
Xfanout388 _04945_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_8
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _03712_ net341 net338 _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_107_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _03437_ net341 net338 _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__o211a_4
XANTENNA__09684__A1 _03462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11710_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12690_ clknet_leaf_50_clk _00254_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07695__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11352__B top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ _05479_ _05505_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07447__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ _05399_ _05405_ _05438_ _05403_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a22o_2
XFILLER_0_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ clknet_leaf_115_clk _00875_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ net2083 net231 net362 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__mux2_1
XANTENNA__10683__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13242_ clknet_leaf_18_clk _00806_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10454_ net244 net2075 net372 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13173_ clknet_leaf_5_clk _00737_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10385_ net256 net1824 net327 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12124_ _05981_ _05990_ _05992_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__and3b_1
XANTENNA__06973__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _05903_ _05905_ _05922_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__nor3_1
X_11006_ net1201 _05019_ net535 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__mux2_1
XANTENNA__06725__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10858__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ clknet_leaf_103_clk _00521_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09675__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11908_ _05740_ _05758_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07686__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ clknet_leaf_110_clk _00452_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__A1 top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ _05673_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12731__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ clknet_leaf_119_clk _01073_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10593__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10993__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07030_ top.DUT.register\[21\]\[11\] net574 net601 top.DUT.register\[10\]\[11\] _02156_
+ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a221o_1
XFILLER_0_180_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08981_ _03146_ net592 net1233 net868 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06964__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ top.DUT.register\[9\]\[16\] net630 net616 top.DUT.register\[30\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_149_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07863_ net808 net493 net463 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__o21a_2
XANTENNA__06716__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06814_ top.DUT.register\[31\]\[24\] net784 net542 top.DUT.register\[22\]\[24\] _01940_
+ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a221o_1
X_09602_ top.a1.state\[1\] net893 top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04634_
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07794_ _02914_ _02916_ _02918_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_162_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ _04552_ _04553_ _04551_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06745_ top.DUT.register\[22\]\[25\] net752 net713 top.DUT.register\[30\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout260_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _04502_ _04503_ _04501_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06676_ top.DUT.register\[14\]\[27\] net611 net599 top.DUT.register\[10\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a22o_1
XANTENNA__08874__C1 _03970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07141__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ _03320_ _03324_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_35_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09395_ top.pc\[20\] _04425_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__nand2_1
XANTENNA__07429__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ net303 _03294_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ _03399_ _03400_ net301 vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07228_ top.DUT.register\[16\]\[15\] net635 net599 top.DUT.register\[10\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ top.DUT.register\[27\]\[13\] net777 net757 top.DUT.register\[11\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10170_ net256 net2305 net409 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
XANTENNA__07601__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10803__Y _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06955__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13607__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1109 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_2
Xfanout130 _05714_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout141 net143 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_2
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
Xfanout163 _04879_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 _04850_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_1
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06707__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 net198 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
X_13860_ net1151 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12811_ clknet_leaf_32_clk _00375_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10678__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ clknet_leaf_67_clk _01334_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07668__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12742_ clknet_leaf_9_clk _00306_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07132__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12673_ clknet_leaf_24_clk _00237_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11624_ _05462_ _05492_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08672__A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11555_ _05413_ _05415_ _05419_ _05421_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_42_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09290__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10506_ net168 net2232 net365 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__mux2_1
XANTENNA__07840__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11486_ _05301_ _05333_ _05306_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_52_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13225_ clknet_leaf_12_clk _00789_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ net184 top.DUT.register\[16\]\[22\] net326 vssd1 vssd1 vccd1 vccd1 _00624_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07199__A2 _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12192__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ clknet_leaf_41_clk _00720_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ net1777 net142 net394 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06946__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12107_ _05951_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13087_ clknet_leaf_114_clk _00651_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10299_ net2213 net146 net402 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
XANTENNA__07776__A_N net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__X _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ _05888_ _05890_ _05896_ _05901_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__or4_1
XANTENNA__12430__Q top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07371__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06530_ net900 _01573_ _01590_ net801 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__and4b_4
XFILLER_0_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07123__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06461_ top.a1.instruction\[3\] net834 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08871__A2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08200_ _03322_ _03325_ net278 vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09180_ _04235_ _04236_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__xnor2_1
X_06392_ _01498_ net791 _01505_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__and3_4
XFILLER_0_172_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ _03156_ _03160_ _03154_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or3b_1
XANTENNA__08623__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ _03186_ net273 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__nor2_1
XANTENNA__06306__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07013_ top.DUT.register\[25\]\[11\] net773 net682 top.DUT.register\[7\]\[11\] _02137_
+ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09584__B1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06937__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ net1276 net870 _02398_ net594 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__a22o_1
X_07915_ top.DUT.register\[25\]\[16\] net772 net684 top.DUT.register\[7\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a22o_1
X_08895_ net475 _03979_ _03992_ net472 vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__o22ai_1
XANTENNA_fanout475_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ top.DUT.register\[24\]\[18\] net551 net602 top.DUT.register\[10\]\[18\] _02972_
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a221o_1
XANTENNA__07898__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07362__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09639__A1 top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _02255_ _02274_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout642_A _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06570__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06728_ _01847_ _01849_ _01851_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__or4_1
X_09516_ _04535_ _04536_ _04537_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ _04486_ _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09859__Y _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06659_ top.DUT.register\[31\]\[27\] net743 net735 top.DUT.register\[24\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout907_A top.i_ready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09378_ top.a1.instruction\[31\] _01615_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08329_ _03450_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11340_ top.a1.dataIn\[19\] _05204_ _05206_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11271_ top.a1.row1\[123\] _05106_ _05108_ top.a1.row1\[11\] _05147_ vssd1 vssd1
+ vccd1 vccd1 _05148_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_115_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13010_ clknet_leaf_48_clk _00574_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10222_ net188 net1962 net407 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__mux2_1
X_10153_ net191 net2205 net415 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10084_ net205 net1790 net419 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
XANTENNA_input36_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 top.a1.dataInTemp\[3\] vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07889__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07353__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ net1144 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_202_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06561__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11093__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13774_ clknet_leaf_65_clk _01317_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10986_ top.a1.dataInTemp\[4\] top.a1.data\[0\] net799 vssd1 vssd1 vccd1 vccd1 _05006_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12725_ clknet_leaf_4_clk _00289_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08853__A2 _03949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ clknet_leaf_0_clk _00220_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11607_ _05415_ _05443_ _05463_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a2bb2o_1
X_12587_ clknet_leaf_29_clk _00151_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07813__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11538_ net250 vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold408 top.DUT.register\[4\]\[2\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12425__Q top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold419 top.DUT.register\[28\]\[7\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _05308_ _05319_ net267 vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__and3_1
XANTENNA__10871__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08369__B2 _03490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ clknet_leaf_111_clk _00772_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06650__A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06919__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ clknet_leaf_5_clk _00703_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 top.DUT.register\[3\]\[18\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 top.DUT.register\[5\]\[19\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ top.DUT.register\[20\]\[0\] net747 net720 top.DUT.register\[14\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__a22o_1
XANTENNA__09869__B2 top.a1.dataIn\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ _03386_ _03542_ _03604_ net271 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__o22a_1
XANTENNA__11140__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ net808 _02757_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_179_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06552__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10111__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _02638_ _02686_ _02206_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
XANTENNA__08864__X _03963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ _04328_ _04332_ _04330_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__o21a_1
X_06513_ _01591_ _01626_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__nand2_2
XFILLER_0_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07493_ top.DUT.register\[11\]\[5\] net639 net607 top.DUT.register\[12\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09232_ _02184_ _02212_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06444_ net904 _01569_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09163_ _04219_ _04220_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06375_ _01497_ _01498_ net792 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_157_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ _03239_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_211_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ _02789_ _02830_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__nor2_1
XANTENNA__07804__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08045_ _01569_ _03154_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__and2_2
XANTENNA__10781__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07927__Y _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold920 top.DUT.register\[25\]\[21\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold931 top.DUT.register\[6\]\[23\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold942 top.ramload\[1\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 top.DUT.register\[21\]\[30\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__A2 _03386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold964 top.DUT.register\[24\]\[29\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 top.DUT.register\[29\]\[16\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 top.DUT.register\[5\]\[25\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 top.DUT.register\[25\]\[23\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ net464 _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net866 _01483_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nor2_4
XANTENNA__06791__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ net886 top.pc\[28\] net537 _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a22o_1
XANTENNA__07335__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07829_ top.DUT.register\[16\]\[18\] _01514_ net745 top.DUT.register\[31\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10840_ net1766 net255 net349 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__mux2_1
XANTENNA__10021__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ net1989 net150 net445 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__mux2_1
XANTENNA__08934__B _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ clknet_leaf_61_clk _00077_ net1099 vssd1 vssd1 vccd1 vccd1 top.ramstore\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06846__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13490_ clknet_leaf_48_clk _01054_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06735__A _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12441_ clknet_leaf_94_clk top.ru.next_FetchedData\[25\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[25\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_117_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ net2107 net912 net36 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11323_ _05183_ _05192_ _05186_ _05190_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or4b_2
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10691__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ top.a1.row2\[1\] _05111_ _05119_ top.a1.row1\[17\] _05132_ vssd1 vssd1 vccd1
+ vccd1 _05133_ sky130_fd_sc_hd__a221o_1
X_10205_ net253 net2004 net408 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11185_ net851 _05066_ net531 vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__and3_1
XANTENNA__08771__A1 _03537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07574__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ _04699_ top.DUT.register\[8\]\[3\] net413 vssd1 vssd1 vccd1 vccd1 _00349_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input39_X net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ net262 net2062 net417 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07326__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__A1 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__A3 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_5__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ clknet_leaf_67_clk _01367_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13757_ clknet_leaf_71_clk _01300_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10866__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10969_ top.a1.halfData\[0\] _04991_ _04992_ net844 vssd1 vssd1 vccd1 vccd1 _04993_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12708_ clknet_leaf_39_clk _00272_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ clknet_leaf_73_clk _01236_ net1090 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__B1 _03164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12639_ clknet_leaf_111_clk _00203_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09787__B1 _04407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06160_ top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 top.DUT.register\[11\]\[9\] vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 top.ramaddr\[2\] vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 top.DUT.register\[14\]\[24\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 top.a1.row1\[112\] vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 top.DUT.register\[14\]\[14\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11346__B1 top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout707 _01533_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10106__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ net802 _04847_ _04848_ _04843_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__a31o_1
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
Xfanout729 net730 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_8
X_08801_ _03265_ _03285_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__nand2_1
X_09781_ net215 top.DUT.register\[1\]\[17\] net437 vssd1 vssd1 vccd1 vccd1 _00139_
+ sky130_fd_sc_hd__mux2_1
X_06993_ net512 _02118_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__and2_1
XANTENNA__11148__D _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08732_ _02079_ net468 _03484_ _03771_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o22a_1
XANTENNA__07317__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09711__B1 _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _03350_ _03770_ _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08100__A _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08959__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07614_ top.DUT.register\[3\]\[2\] net785 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__and2_1
X_08594_ _02275_ _02319_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ top.DUT.register\[25\]\[4\] net773 net683 top.DUT.register\[7\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XANTENNA__10776__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08817__A2 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout438_A _04681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07476_ top.DUT.register\[6\]\[5\] net763 net671 top.DUT.register\[16\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06427_ net790 _01503_ _01506_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__and3_4
X_09215_ _04262_ _04265_ _04263_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout605_A _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09778__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _04192_ _04195_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a21oi_1
X_06358_ top.lcd.cnt_500hz\[13\] _01487_ top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1
+ vccd1 top.lcd.lcd_en sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ _01909_ _02879_ net468 _03415_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or4b_1
X_06289_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_112_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ _01480_ _01581_ _01607_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_96_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 top.DUT.register\[25\]\[9\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 top.DUT.register\[27\]\[4\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold772 top.DUT.register\[19\]\[24\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold783 top.DUT.register\[26\]\[7\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10016__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 top.a1.row1\[15\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ net2036 net217 net429 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA__06764__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ clknet_leaf_14_clk _00554_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09702__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11941_ _05809_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__nand2_2
X_11872_ _05705_ net131 vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13611_ clknet_leaf_98_clk net1176 net981 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10686__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ net1563 net205 net355 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_118_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ clknet_leaf_24_clk _01106_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ net180 net1775 net374 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ net223 net1926 net377 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
X_13473_ clknet_leaf_28_clk _01037_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ clknet_leaf_100_clk top.ru.next_FetchedData\[8\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[8\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09776__A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12355_ top.pad.button_control.r_counter\[11\] _06141_ vssd1 vssd1 vccd1 vccd1 _06142_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07795__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ top.a1.row1\[63\] _05112_ _05169_ _05175_ _05178_ vssd1 vssd1 vccd1 vccd1
+ _05179_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_39_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12286_ _01436_ net588 _06099_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__and3_1
XANTENNA__11328__B1 top.a1.dataIn\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11237_ _05092_ _05110_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_52_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ top.a1.dataInTemp\[6\] top.a1.data\[6\] net799 vssd1 vssd1 vccd1 vccd1 _05072_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output67_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06755__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ net1524 net187 net460 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
X_11099_ net71 net859 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09016__A _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07180__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ clknet_leaf_68_clk _01352_ net1104 vssd1 vssd1 vccd1 vccd1 top.pad.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10596__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_109_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10067__A0 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07330_ top.DUT.register\[11\]\[8\] net755 net712 top.DUT.register\[30\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11712__C top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07483__A1 top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07261_ top.DUT.register\[7\]\[14\] net554 net550 top.DUT.register\[24\]\[14\] _02387_
+ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a221o_1
X_09000_ _03979_ _03998_ _04017_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__and4_1
XANTENNA__12909__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06212_ top.ru.state\[6\] top.busy_o top.ru.state\[3\] vssd1 vssd1 vccd1 vccd1 _01428_
+ sky130_fd_sc_hd__a21o_2
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_154_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07192_ _02298_ _02317_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07786__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ net835 _04585_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07538__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
XANTENNA__12497__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09833_ net834 _04485_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__o21bai_1
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
Xfanout548 _01661_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_4
Xfanout559 _01653_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_4
XANTENNA__06746__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Right_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_206_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout388_A _04945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06210__A2 top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _04769_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__or2_1
X_06976_ top.DUT.register\[16\]\[20\] net638 net617 top.DUT.register\[30\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a22o_1
X_08715_ _03208_ _03213_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__nand2_1
X_09695_ net245 net2176 net440 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08646_ _03755_ _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__or2_2
XFILLER_0_194_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07710__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout722_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ net1271 net839 net817 _03690_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07528_ top.DUT.register\[31\]\[4\] net783 net622 top.DUT.register\[26\]\[4\] _02654_
+ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12146__A_N top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07459_ _02567_ _02585_ net806 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_2
XANTENNA__11270__A2 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ net183 net1953 net371 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
X_09129_ _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ _05989_ _06003_ _05997_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_94_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06985__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ _05939_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nand2_1
Xhold580 top.DUT.register\[31\]\[28\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07529__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold591 top.DUT.register\[11\]\[1\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ net32 net831 net830 net1829 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__a22o_1
XANTENNA__07844__A _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__B _03768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_204_Left_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12973_ clknet_leaf_23_clk _00537_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11924_ _05775_ _05791_ _05793_ _05773_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07162__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11855_ _05687_ net130 vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ net1411 net260 net353 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__mux2_1
XANTENNA__06195__A top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11786_ _05629_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08961__A1_N net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13525_ clknet_leaf_5_clk _01089_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10737_ net144 net1716 net382 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__mux2_1
XANTENNA__08662__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08681__Y _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13456_ clknet_leaf_121_clk _01020_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08614__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10668_ net1946 net169 net451 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__mux2_1
X_12407_ clknet_leaf_81_clk _00043_ net1013 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12210__A1 top.a1.row2\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10599_ net192 net2069 net388 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
X_13387_ clknet_leaf_29_clk _00951_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XANTENNA__08965__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12338_ _06130_ _06131_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__nor2_1
XANTENNA__06976__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__Q top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ net1213 _06087_ _06089_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06830_ top.DUT.register\[28\]\[23\] net651 net643 top.DUT.register\[17\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire523_A _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07940__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ top.DUT.register\[16\]\[25\] net636 net612 top.DUT.register\[14\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a22o_1
X_08500_ net888 top.pc\[10\] net537 _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__a22o_1
X_09480_ net517 _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__nand2b_1
X_06692_ _01818_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__inv_2
XANTENNA__07153__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08431_ net479 _03534_ _03550_ net476 _03547_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06900__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ net311 _03483_ _03467_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_148_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08248__A3 _03127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07313_ top.DUT.register\[27\]\[9\] net596 net541 top.DUT.register\[22\]\[9\] _02439_
+ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08293_ _03416_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07244_ _02368_ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06392__X _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07175_ top.DUT.register\[21\]\[13\] net574 net650 top.DUT.register\[13\]\[13\] _02301_
+ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12201__B2 top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__B2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06967__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__A3 _03537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12607__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06431__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A_N _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _02760_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_167_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 _02711_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_4
Xfanout323 _04957_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_8
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _04964_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_8
Xfanout356 _04962_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_4
X_09816_ net834 _04452_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__o21bai_1
Xfanout367 _04959_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 _04949_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_4
XFILLER_0_185_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout389 _04944_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_6
XFILLER_0_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07931__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ net802 _04754_ _04755_ _04750_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a31o_1
X_06959_ top.DUT.register\[9\]\[20\] net710 net669 top.DUT.register\[5\]\[20\] _02085_
+ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout937_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_190_Right_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ top.pc\[3\] net803 net343 _04697_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a211o_1
XANTENNA__09684__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08629_ net474 _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nor2_1
XANTENNA__08892__B1 _03989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11640_ _05478_ _05505_ _05475_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_194_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _05425_ _05433_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a21o_2
XFILLER_0_147_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ clknet_leaf_14_clk _00874_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10522_ net1682 net237 net361 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13241_ clknet_leaf_35_clk _00805_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ net247 net1792 net369 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13172_ clknet_leaf_60_clk _00736_ net1102 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10384_ net261 net1852 net327 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__mux2_1
XANTENNA__06958__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12123_ _05990_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__and2_1
X_12054_ _05905_ _05922_ _05903_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21a_1
XANTENNA__08713__A2_N net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ top.a1.dataIn\[10\] net848 net843 _05018_ vssd1 vssd1 vccd1 vccd1 _05019_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10204__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout890 top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07922__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06477__X _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12956_ clknet_leaf_55_clk _00520_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07135__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11907_ _05757_ _05759_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ clknet_leaf_105_clk _00451_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10690__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11838_ _05658_ _05662_ _05677_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12428__Q top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10874__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__C1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _05603_ _05620_ _05637_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_40_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13508_ clknet_leaf_43_clk _01072_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07749__A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08344__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10993__A1 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13439_ clknet_leaf_114_clk _01003_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06661__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12195__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06949__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12700__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ net1309 net868 _01689_ net594 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07931_ top.DUT.register\[24\]\[16\] net549 net612 top.DUT.register\[14\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_149_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07862_ _02973_ _02986_ _02987_ _02988_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__nor4_1
XANTENNA__10114__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07374__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__inv_2
X_06813_ top.DUT.register\[19\]\[24\] net634 net780 top.DUT.register\[15\]\[24\] _01931_
+ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a221o_1
X_07793_ top.DUT.register\[9\]\[19\] net709 net676 top.DUT.register\[18\]\[19\] _02919_
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06744_ top.DUT.register\[29\]\[25\] net701 _01869_ _01870_ vssd1 vssd1 vccd1 vccd1
+ _01871_ sky130_fd_sc_hd__a211o_1
XANTENNA__06387__X _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09463_ top.pc\[24\] _04493_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__or2_1
X_06675_ top.DUT.register\[28\]\[27\] net651 net639 top.DUT.register\[11\]\[27\] _01801_
+ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout253_A _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08414_ net317 _03533_ _03530_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09394_ _04418_ _04420_ _04417_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_35_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08345_ net285 _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10784__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_31_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ _03309_ _03322_ net281 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
XANTENNA__12859__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10984__A1 top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10984__B2 _05004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06652__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ top.DUT.register\[20\]\[15\] net576 net567 top.DUT.register\[4\]\[15\] _02353_
+ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ top.DUT.register\[8\]\[13\] net742 net737 top.DUT.register\[24\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout887_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07089_ top.DUT.register\[8\]\[10\] net568 net541 top.DUT.register\[22\]\[10\] _02215_
+ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a221o_1
Xfanout1107 net1109 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_196_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout131 _05714_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_98_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09354__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12777__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout153 net155 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10024__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout164 _04868_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07365__A0 _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout175 net178 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_2
Xfanout186 _04831_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07681__X _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_137_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12810_ clknet_leaf_40_clk _00374_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13790_ clknet_leaf_67_clk _01333_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06297__X _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__B1 _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ clknet_leaf_118_clk _00305_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12672_ clknet_leaf_45_clk _00236_ net1080 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11623_ _05462_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__or2_1
XANTENNA__06891__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10694__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08617__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire510 _02161_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_2
X_11554_ _05413_ _05415_ _05419_ _05421_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_146_Left_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10975__A1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12529__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10505_ net172 net2275 net367 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__mux2_1
XANTENNA__06643__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11485_ _05306_ _05333_ _05301_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_133_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ clknet_leaf_35_clk _00788_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10436_ net189 net1764 net326 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09593__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ clknet_leaf_41_clk _00719_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09593__B2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10367_ net1723 net144 net396 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12106_ top.a1.dataIn\[3\] _05961_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_209_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13086_ clknet_leaf_14_clk _00650_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10298_ net1583 net153 net403 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_89_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12037_ _05888_ _05901_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__or2_1
XANTENNA__09008__B _03843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_155_Left_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07356__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__B2 top.busy_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07751__B _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ clknet_leaf_29_clk _00503_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06367__B net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06460_ top.a1.instruction\[3\] net834 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06882__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06391_ _01497_ net792 _01508_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__and3_4
XANTENNA__11207__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_164_Left_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08130_ _03175_ _03154_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__and2b_2
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ net322 net310 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__nand2_1
XANTENNA__06634__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ top.DUT.register\[12\]\[11\] net583 net673 top.DUT.register\[16\]\[11\] _02138_
+ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07485__Y _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11391__A1 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07595__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ net523 net591 net1210 net870 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08103__A _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_173_Left_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09336__B2 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ top.DUT.register\[4\]\[16\] net770 _01520_ top.DUT.register\[17\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__a22o_1
XANTENNA__07347__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ _03104_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__nand2_1
X_13846__1147 vssd1 vssd1 vccd1 vccd1 net1147 _13846__1147/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ top.DUT.register\[1\]\[18\] net658 net618 top.DUT.register\[30\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a22o_1
XANTENNA__10779__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A _04958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__C _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11464__A top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A _03339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07776_ net503 _02447_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_88_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09515_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__nand2_1
X_06727_ top.DUT.register\[29\]\[26\] net665 net625 top.DUT.register\[25\]\[26\] _01853_
+ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout635_A _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09446_ top.pc\[23\] _04476_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_182_Left_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06845__X _01972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06658_ top.DUT.register\[28\]\[27\] net584 net708 top.DUT.register\[9\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12295__A _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06873__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ _02971_ _04407_ _04410_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout802_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06589_ top.DUT.register\[2\]\[29\] net662 net649 top.DUT.register\[13\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08328_ _02685_ _03413_ _03419_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nand3_1
XFILLER_0_191_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06625__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _03224_ _03226_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__nand2_1
XANTENNA__10019__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11270_ net885 _05103_ _05112_ top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 _05147_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10221_ net192 net2143 net408 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__mux2_1
XANTENNA__07586__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ net205 net2244 net416 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
XANTENNA__07050__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10083_ net212 net1609 net420 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__mux2_1
XANTENNA__08948__A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 top.a1.dataInTemp\[0\] vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07889__A1 top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ net1111 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_202_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13773_ clknet_leaf_65_clk _01316_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10985_ net2238 _05005_ net535 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12724_ clknet_leaf_60_clk _00288_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09779__A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ clknet_leaf_18_clk _00219_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11606_ _05413_ _05415_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__nand2_1
X_12586_ clknet_leaf_38_clk _00150_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06616__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11537_ _05399_ _05405_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12942__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold409 top.DUT.register\[18\]\[31\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
X_11468_ top.a1.dataIn\[15\] _05334_ _05335_ _05336_ vssd1 vssd1 vccd1 vccd1 _05338_
+ sky130_fd_sc_hd__o211a_1
Xmax_cap128 _05862_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_1
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ clknet_leaf_107_clk _00771_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ net254 net1991 net325 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__mux2_1
XANTENNA__09566__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ _05236_ _05237_ _05256_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07577__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13138_ clknet_leaf_49_clk _00702_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07041__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13069_ clknet_leaf_25_clk _00633_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07329__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1109 top.DUT.register\[18\]\[0\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_146_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09869__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__A2 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ _02743_ _02754_ _02755_ _02756_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_179_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07561_ _02687_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__inv_2
X_09300_ _02380_ _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__xor2_1
X_06512_ _01573_ _01631_ _01634_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__and3_4
X_07492_ top.DUT.register\[2\]\[5\] net659 net651 top.DUT.register\[28\]\[5\] _02618_
+ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_192_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ _04283_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__xnor2_1
X_06443_ net905 _01476_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__nand2_2
XFILLER_0_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06374_ top.a1.instruction\[19\] net810 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nand2_1
X_09162_ _04220_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08113_ _02339_ net290 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11061__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09093_ _02835_ _02876_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_211_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout216_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ _03169_ _03170_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__and2_1
XANTENNA__07280__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold910 top.DUT.register\[11\]\[8\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold921 top.DUT.register\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 top.DUT.register\[28\]\[5\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 top.DUT.register\[21\]\[1\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 top.DUT.register\[31\]\[13\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 top.DUT.register\[31\]\[12\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 top.DUT.register\[29\]\[0\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold998 top.DUT.register\[19\]\[12\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _04685_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout585_A _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08780__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net1263 net1163 _04040_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11116__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08877_ _03974_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ top.DUT.register\[20\]\[18\] net750 net734 top.DUT.register\[19\]\[18\] _02952_
+ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_86_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_190_Left_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07759_ _02885_ _02685_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__Y _03878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10627__A0 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07099__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10770_ net143 net2019 net375 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09493__B1 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09429_ _04455_ _04457_ _04454_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06846__A2 _01972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__B _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ clknet_leaf_94_clk top.ru.next_FetchedData\[24\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08054__A1_N _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09796__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__A2 _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net2182 net912 net35 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11322_ top.a1.dataIn\[23\] _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09548__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ net891 top.a1.row1\[113\] _05105_ _05129_ vssd1 vssd1 vccd1 vccd1 _05132_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06470__B top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__C1 _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ net255 net1691 net405 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__mux2_1
XANTENNA__07023__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08220__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _01409_ _04977_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__or2_2
XFILLER_0_207_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08771__A2 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ net259 top.DUT.register\[8\]\[2\] net413 vssd1 vssd1 vccd1 vccd1 _00348_
+ sky130_fd_sc_hd__mux2_1
X_10066_ net264 net1476 net419 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08523__A2 _03619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07731__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13825_ clknet_leaf_67_clk _01366_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08684__Y _03793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13756_ clknet_leaf_73_clk _01299_ net1094 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10968_ top.a1.dataInTemp\[0\] net800 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12707_ clknet_leaf_33_clk _00271_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12544__RESET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13687_ clknet_leaf_73_clk _01235_ net1094 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ net2318 net154 net347 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08039__A1 _03127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ clknet_leaf_15_clk _00202_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13845__1146 vssd1 vssd1 vccd1 vccd1 net1146 _13845__1146/LO sky130_fd_sc_hd__conb_1
XFILLER_0_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06364__C net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ clknet_leaf_37_clk _00133_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07798__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold206 top.DUT.register\[14\]\[12\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 top.DUT.register\[23\]\[13\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 top.DUT.register\[24\]\[8\] vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 top.DUT.register\[11\]\[20\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout708 net711 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout719 _01529_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
X_08800_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__inv_2
X_09780_ _03776_ net342 net339 _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ net512 _02118_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__nor2_1
X_08731_ _02078_ net485 net487 _02077_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10122__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ _03034_ net485 net470 _03035_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07722__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ top.DUT.register\[21\]\[2\] net572 net623 top.DUT.register\[25\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ net482 _03705_ _03699_ _03697_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__o211a_1
XANTENNA__08594__Y _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout166_A _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07544_ top.DUT.register\[28\]\[4\] net586 net582 top.DUT.register\[12\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
XANTENNA__08278__B2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06395__X _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09475__B1 _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08483__A2_N _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06828__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07475_ top.DUT.register\[23\]\[5\] net696 _02596_ _02601_ vssd1 vssd1 vccd1 vccd1
+ _02602_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_81_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1075_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09214_ top.pc\[9\] _04254_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__xnor2_1
X_06426_ _01496_ net793 _01505_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09145_ _02641_ _02682_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__xor2_1
X_06357_ _01485_ _01486_ top.lcd.cnt_500hz\[11\] top.lcd.cnt_500hz\[12\] vssd1 vssd1
+ vccd1 vccd1 _01487_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_20_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09778__B2 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07789__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06288_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 _01436_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08450__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09076_ _01821_ _01865_ _02589_ _03525_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__or4bb_1
XANTENNA__08450__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08027_ _01607_ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_96_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11189__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 top.DUT.register\[23\]\[26\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 top.DUT.register\[17\]\[3\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 top.DUT.register\[17\]\[29\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold773 top.DUT.register\[9\]\[21\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08202__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 top.DUT.register\[19\]\[0\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 top.DUT.register\[13\]\[11\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ net1430 net229 net430 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
X_08929_ net487 _03742_ _04024_ _03151_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09702__A1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _05774_ _05787_ _05789_ _05767_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__or4b_1
XANTENNA__10032__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07713__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _05703_ _05740_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_196_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ clknet_leaf_98_clk net1255 net981 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10822_ net2185 net213 net356 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09122__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ clknet_leaf_119_clk _01105_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13640__Q net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06819__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10753_ net196 net1465 net375 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13472_ clknet_leaf_49_clk _01036_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07492__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13143__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ net231 net1974 net378 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ clknet_leaf_97_clk top.ru.next_FetchedData\[7\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_164_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12354_ _06141_ net796 _06140_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__and3b_1
XANTENNA__08441__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11305_ _05093_ _05176_ _05177_ net881 _05166_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10207__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12285_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 _06099_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09792__A top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ net891 net880 _05114_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net1289 net533 net525 _05071_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__a22o_1
X_10118_ net1355 net192 net461 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
X_11098_ net917 net2033 net852 _05035_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10049_ net213 net2323 net423 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10877__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13808_ clknet_leaf_68_clk _01351_ net1104 vssd1 vssd1 vccd1 vccd1 top.pad.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09457__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ clknet_leaf_74_clk _01282_ net1018 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11712__D top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07260_ top.DUT.register\[12\]\[14\] net609 net597 top.DUT.register\[27\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a22o_1
XANTENNA__08680__A1 _03386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06211_ net34 _01427_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07191_ _02298_ _02317_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_154_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__A1 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10117__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09901_ _04881_ _04885_ _04893_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__nand3_1
XFILLER_0_111_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12660__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload20_A clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _04493_ net526 net332 top.a1.dataIn\[23\] net335 vssd1 vssd1 vccd1 vccd1
+ _04832_ sky130_fd_sc_hd__a221o_1
Xfanout527 _04745_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
Xfanout549 _01661_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07943__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09207__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ top.pc\[16\] _04379_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__nor2_1
XANTENNA__08111__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ top.DUT.register\[4\]\[20\] net565 net626 top.DUT.register\[25\]\[20\] _02101_
+ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout283_A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08714_ _02121_ net470 _03446_ _03770_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a221o_1
XANTENNA__11098__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09694_ _03521_ net340 net336 _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__o211a_2
XFILLER_0_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08645_ _03075_ net486 net522 _03752_ _03740_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout450_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10787__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ net889 top.pc\[13\] net537 _03689_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06566__A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07527_ top.DUT.register\[19\]\[4\] net633 net780 top.DUT.register\[15\]\[4\] _02644_
+ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a221o_1
XANTENNA__11191__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout715_A _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ _02580_ _02582_ _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__or3_2
XFILLER_0_162_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07474__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06409_ net792 _01503_ _01508_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_98_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09596__B top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07389_ _02507_ _02515_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__nor2_8
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09128_ top.pc\[3\] _02739_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and2_1
XANTENNA__07226__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09883__Y _04879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09059_ _04120_ _03149_ _02587_ net485 vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__and4b_1
XFILLER_0_130_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07684__X _02811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12070_ _05919_ _05931_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__xnor2_1
Xhold570 top.DUT.register\[8\]\[21\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 top.DUT.register\[27\]\[16\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08499__Y _03616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 top.DUT.register\[13\]\[2\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net31 net841 net811 net1415 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__o22a_1
XANTENNA__09923__A1 _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__A2 top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13844__1145 vssd1 vssd1 vccd1 vccd1 net1145 _13844__1145/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_125_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ clknet_leaf_9_clk _00536_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09687__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11923_ _05772_ _05791_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10697__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11854_ _05722_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10805_ net2166 net263 net355 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
X_11785_ _05626_ _05638_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_171_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13524_ clknet_leaf_47_clk _01088_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ net153 net1765 net384 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07465__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06673__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13455_ clknet_leaf_51_clk _01019_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10667_ net1384 net173 net451 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12406_ clknet_leaf_81_clk _00042_ net1006 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08414__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07217__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13386_ clknet_leaf_34_clk _00950_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12210__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10598_ net203 net1690 net388 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12337_ net1854 _06128_ net795 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__o21ai_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__08958__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ net1213 _06087_ net1108 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ net879 top.lcd.nextState\[4\] _05095_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__and3_1
XANTENNA_max_cap513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ _05984_ _04976_ net845 net2082 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__a2bb2o_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__07925__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09027__A _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06760_ top.DUT.register\[11\]\[25\] net640 net557 top.DUT.register\[6\]\[25\] _01886_
+ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a221o_1
XANTENNA__09678__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06691_ _01797_ _01816_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__and2_2
XFILLER_0_203_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_201_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__nand2_1
XANTENNA__10400__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08361_ net303 _03348_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07312_ top.DUT.register\[17\]\[9\] net644 net627 top.DUT.register\[9\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07456__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ _02884_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08805__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06664__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07243_ top.DUT.register\[6\]\[14\] net765 net730 top.DUT.register\[10\]\[14\] _02369_
+ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07208__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ top.DUT.register\[16\]\[13\] net638 net601 top.DUT.register\[10\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1038_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_7__f_clk_X clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net318 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
Xfanout324 _04957_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
Xfanout335 _04717_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
Xfanout346 _04964_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07916__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _04460_ net526 net332 top.a1.dataIn\[21\] net334 vssd1 vssd1 vccd1 vccd1
+ _04817_ sky130_fd_sc_hd__a221o_1
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 net360 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_6
Xfanout368 _04959_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_4
Xfanout379 _04949_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_6
XANTENNA_fanout665_A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ _04740_ _04742_ _04753_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__o21bai_1
X_06958_ top.DUT.register\[25\]\[20\] net773 net750 top.DUT.register\[20\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09677_ _01568_ _04182_ _04183_ net794 top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1
+ _04697_ sky130_fd_sc_hd__a32o_1
X_06889_ top.DUT.register\[2\]\[22\] net661 net598 top.DUT.register\[27\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10310__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ _03737_ _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06296__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07695__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__B2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ _02320_ _03672_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ _05439_ _05436_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08644__A1 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13435__RESET_B net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06655__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ net1541 net240 net361 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13240_ clknet_leaf_108_clk _00804_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ net251 net1903 net371 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06407__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ clknet_leaf_1_clk _00735_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10383_ net264 net1689 net329 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12122_ _05976_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12053_ _05905_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ top.a1.data\[6\] top.a1.dataInTemp\[10\] net797 vssd1 vssd1 vccd1 vccd1 _05018_
+ sky130_fd_sc_hd__mux2_1
Xfanout880 top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_2
Xfanout891 top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_2
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input14_X net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ clknet_leaf_58_clk _00519_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11906_ _05770_ _05771_ _05773_ _05767_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__or4b_4
XFILLER_0_197_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10220__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07686__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ clknet_leaf_2_clk _00450_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06894__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ _05663_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_138_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _05614_ _05635_ _05636_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__a21o_2
XFILLER_0_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13507_ clknet_leaf_50_clk _01071_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10719_ net207 net2257 net381 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ _05540_ _05546_ _05551_ _05559_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__nand4_1
XFILLER_0_126_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10993__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13438_ clknet_leaf_14_clk _01002_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12444__Q top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10890__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ clknet_leaf_37_clk _00933_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06949__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ top.DUT.register\[2\]\[16\] net660 net557 top.DUT.register\[6\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ top.DUT.register\[2\]\[18\] net662 net570 top.DUT.register\[8\]\[18\] _02974_
+ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__a221o_1
XANTENNA__12579__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ top.a1.state\[2\] _04628_ net893 top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04632_ sky130_fd_sc_hd__or4bb_1
X_06812_ top.DUT.register\[6\]\[24\] net558 net602 top.DUT.register\[10\]\[24\] _01938_
+ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ top.DUT.register\[22\]\[19\] net754 net679 top.DUT.register\[13\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ top.pc\[27\] _04532_ top.pc\[28\] vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__a21oi_1
X_06743_ top.DUT.register\[6\]\[25\] net764 net674 top.DUT.register\[18\]\[25\] _01866_
+ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09462_ top.pc\[24\] _04493_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__nand2_1
X_06674_ top.DUT.register\[17\]\[27\] net643 net615 top.DUT.register\[30\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a22o_1
XANTENNA__08874__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08413_ net311 net299 _03429_ _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_195_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06885__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09393_ net136 _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11750__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08344_ _03271_ _03287_ net298 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07429__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06637__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ _03315_ _03325_ net288 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout413_A _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10984__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07226_ top.DUT.register\[2\]\[15\] net659 net651 top.DUT.register\[28\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13843__1144 vssd1 vssd1 vccd1 vccd1 net1144 _13843__1144/LO sky130_fd_sc_hd__conb_1
XFILLER_0_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08929__A2 _03742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ top.DUT.register\[29\]\[13\] net703 net694 top.DUT.register\[21\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09874__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10372__Y _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07601__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ top.DUT.register\[29\]\[10\] net663 net548 top.DUT.register\[24\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout782_A _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11197__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__A_N net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1109 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10305__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout132 net135 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08960__A1_N _02231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 _04915_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
Xfanout165 _04868_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_1
XANTENNA__07365__A1 _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 net178 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 _04820_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
Xfanout198 _04757_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_2
X_09729_ top.pc\[13\] _04329_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09511__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ clknet_leaf_39_clk _00304_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10040__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06876__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12671_ clknet_leaf_114_clk _00235_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11622_ _05474_ _05479_ _05483_ _05467_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a211o_1
XFILLER_0_139_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire500 _02469_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
XFILLER_0_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _05419_ _05421_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__and2_1
XANTENNA__09290__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10975__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ net175 net2243 net365 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07840__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11484_ _05301_ _05333_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13223_ clknet_leaf_27_clk _00787_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10435_ net193 net2234 net326 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07053__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ clknet_leaf_41_clk _00718_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ net1445 net153 net394 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12105_ _05969_ _05970_ _05973_ _05958_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__and4b_4
XFILLER_0_20_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06800__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ clknet_leaf_107_clk _00649_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10215__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10297_ net2050 net159 net403 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
X_12036_ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__inv_2
XANTENNA__09008__C _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12938_ clknet_leaf_38_clk _00502_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10885__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12869_ clknet_leaf_118_clk _00433_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06390_ net793 _01505_ _01506_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__and3_4
XANTENNA__08208__X _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06619__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08060_ net316 net285 vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_190_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07292__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07831__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ top.DUT.register\[4\]\[11\] net768 net733 top.DUT.register\[19\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06670__Y _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07044__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12921__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10125__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ net505 net592 net1161 net870 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_164_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07913_ top.DUT.register\[19\]\[16\] net732 net693 top.DUT.register\[21\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a22o_1
X_08893_ _01736_ _01775_ _03103_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__nand3_1
XANTENNA__08544__B1 _03652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__C1 _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07844_ _02970_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__inv_2
XANTENNA__06398__X _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07775_ _02361_ _02901_ _02897_ _02896_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_88_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout363_A _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06570__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ top.pc\[27\] _04543_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__nand2_1
X_06726_ top.DUT.register\[15\]\[26\] net780 _01841_ _01852_ vssd1 vssd1 vccd1 vccd1
+ _01853_ sky130_fd_sc_hd__a211o_1
X_09445_ top.pc\[23\] _04476_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__nor2_1
X_06657_ top.DUT.register\[4\]\[27\] net767 net720 top.DUT.register\[14\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10795__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout628_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ _04418_ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__xnor2_1
X_06588_ top.DUT.register\[15\]\[29\] _01655_ net783 top.DUT.register\[31\]\[29\]
+ _01714_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a221o_1
X_08327_ _03413_ _03419_ _02685_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08075__A2 _03127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07283__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ net287 _03168_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout997_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07209_ top.DUT.register\[27\]\[15\] net775 net727 top.DUT.register\[10\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a22o_1
X_08189_ _03313_ _03314_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07035__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ net204 net2335 net407 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ net212 net1907 net415 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XANTENNA__10035__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10082_ net215 net2281 net417 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__mux2_1
XANTENNA__07889__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ net72 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13643__Q net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06561__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13772_ clknet_leaf_66_clk _01315_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10984_ top.a1.dataIn\[3\] net848 _05003_ _05004_ _04991_ vssd1 vssd1 vccd1 vccd1
+ _05005_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06849__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12723_ clknet_leaf_1_clk _00287_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07510__A1 top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12654_ clknet_leaf_117_clk _00218_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11605_ _05421_ _05463_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12585_ clknet_leaf_2_clk _00149_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11536_ _05344_ _05402_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07813__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11467_ _05335_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__nand2_1
XANTENNA__07026__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ clknet_leaf_121_clk _00770_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10418_ net257 net1850 net323 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__mux2_1
X_11398_ _05266_ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13137_ clknet_leaf_12_clk _00701_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10349_ net1366 net207 net395 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ clknet_leaf_11_clk _00632_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _05860_ net127 _05861_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10884__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06552__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ top.a1.instruction\[15\] net524 _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08829__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06511_ _01573_ _01631_ _01637_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__and3_4
XFILLER_0_158_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07491_ top.DUT.register\[9\]\[5\] net627 net599 top.DUT.register\[10\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09230_ top.pc\[10\] _02427_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__xnor2_1
X_06442_ net905 _01476_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_83_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _02608_ _02612_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__and2_1
X_06373_ top.a1.instruction\[19\] net810 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08112_ _02380_ net290 vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ _04153_ net534 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_211_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07804__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08043_ net296 net467 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold900 top.DUT.register\[30\]\[27\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold911 top.DUT.register\[27\]\[5\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold922 top.a1.row2\[18\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold933 top.DUT.register\[17\]\[1\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 top.DUT.register\[6\]\[14\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 top.DUT.register\[18\]\[10\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 top.a1.row1\[56\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 top.DUT.register\[2\]\[23\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ top.a1.instruction\[10\] _04675_ top.a1.instruction\[9\] vssd1 vssd1 vccd1
+ vccd1 _04921_ sky130_fd_sc_hd__nand3b_4
XANTENNA_fanout1020_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 top.DUT.register\[22\]\[16\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 top.DUT.register\[5\]\[28\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _04033_ _04037_ _04038_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or4_1
XANTENNA__08401__X _03522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout480_A _03255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06791__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout578_A _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _03938_ _03955_ _03973_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nor3_1
XFILLER_0_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13279__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ top.DUT.register\[8\]\[18\] net742 net688 top.DUT.register\[1\]\[18\] _02953_
+ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A _01518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ _02732_ _02884_ _02733_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__o21ba_1
X_06709_ top.DUT.register\[30\]\[26\] net715 _01826_ _01835_ vssd1 vssd1 vccd1 vccd1
+ _01836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07689_ top.DUT.register\[4\]\[0\] net767 net685 top.DUT.register\[1\]\[0\] _02813_
+ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a221o_1
XANTENNA__09493__B2 _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09428_ _04468_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09359_ top.pc\[18\] _04394_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09819__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07256__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ _01402_ _06151_ net795 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_185_Right_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11321_ top.a1.dataIn\[21\] top.a1.dataIn\[20\] top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 _05191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07008__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11252_ top.a1.row2\[33\] _05107_ _05112_ top.a1.row1\[57\] _05130_ vssd1 vssd1 vccd1
+ vccd1 _05131_ sky130_fd_sc_hd__a221o_1
XANTENNA__08024__A _03127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08756__B1 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ net260 net2333 net405 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__mux2_1
XANTENNA__12542__Q top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__A0 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _01409_ _04977_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ net266 net2149 net416 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10065_ net148 top.DUT.register\[6\]\[0\] net417 vssd1 vssd1 vccd1 vccd1 _00282_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09720__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13824_ clknet_leaf_67_clk _01365_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ net849 net844 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__nor2_1
X_13755_ clknet_leaf_71_clk _01298_ net1094 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_12706_ clknet_leaf_42_clk _00270_ net1077 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07495__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10898_ net1562 net158 net348 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
X_13686_ clknet_leaf_72_clk _01234_ net1095 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_174_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ clknet_leaf_107_clk _00201_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06364__D net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ clknet_leaf_110_clk _00132_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ _05349_ _05363_ _05369_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__or3b_1
XFILLER_0_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12499_ clknet_leaf_81_clk _00066_ net1013 vssd1 vssd1 vccd1 vccd1 top.ramstore\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold207 top.pad.button_control.r_counter\[9\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold218 top.DUT.register\[29\]\[9\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 top.ramstore\[19\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout709 net711 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06222__B2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ net808 net511 net463 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__o21a_1
XANTENNA__06773__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07970__A1 _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ net315 _03470_ _03543_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o21a_1
XANTENNA__10403__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08661_ net321 _03256_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__nand2_4
XANTENNA__09711__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07612_ _01616_ _02737_ _02738_ _02734_ net529 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a32o_4
X_08592_ net320 _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload98_A clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07543_ top.DUT.register\[21\]\[4\] net694 net669 top.DUT.register\[5\]\[4\] _02669_
+ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a221o_1
XANTENNA__09475__B2 top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_A _04890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07486__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07474_ top.DUT.register\[11\]\[5\] net755 net667 top.DUT.register\[5\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09213_ net909 top.pc\[8\] _04268_ net898 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06425_ top.DUT.register\[28\]\[30\] net585 _01538_ _01551_ vssd1 vssd1 vccd1 vccd1
+ _01552_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1068_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _04200_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__xnor2_1
X_06356_ top.lcd.cnt_500hz\[8\] top.lcd.cnt_500hz\[9\] top.lcd.cnt_500hz\[10\] vssd1
+ vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09075_ _03078_ _03171_ _04136_ _02783_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__or4b_1
X_06287_ top.ramload\[31\] net877 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ net903 _01606_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold730 top.ramload\[2\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold741 top.DUT.register\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08738__B1 _03843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout695_A _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold752 top.DUT.register\[8\]\[9\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 top.DUT.register\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold774 top.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap493 _02989_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_2
Xhold785 top.DUT.register\[21\]\[6\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 top.DUT.register\[29\]\[2\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net2138 net180 net430 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
XANTENNA__06764__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net484 net468 _03149_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08859_ _01820_ _01861_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11870_ _05738_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__or2_2
XFILLER_0_211_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ net2063 net218 net353 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_40_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13540_ clknet_leaf_41_clk _01104_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07477__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10752_ net199 net1442 net375 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12537__Q top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13471_ clknet_leaf_114_clk _01035_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10683_ net236 net1388 net377 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12422_ clknet_leaf_97_clk top.ru.next_FetchedData\[6\] net985 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[6\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07229__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08977__B1 _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12353_ top.pad.button_control.r_counter\[10\] top.pad.button_control.r_counter\[9\]
+ _06137_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11304_ net891 _05115_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__nor2_1
X_12284_ top.lcd.cnt_500hz\[0\] net588 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_39_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11235_ net879 top.lcd.nextState\[4\] _05092_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__or3_1
XANTENNA__09792__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07401__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ top.a1.dataInTemp\[5\] top.a1.data\[5\] net799 vssd1 vssd1 vccd1 vccd1 _05071_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net1979 net203 net461 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XANTENNA__10223__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ net70 net857 vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__and2_1
X_10048_ net217 net2052 net421 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__mux2_1
Xhold90 _01321_ vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07180__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ clknet_leaf_64_clk _01350_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_max_cap493_A _02989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11999_ _05811_ _05838_ _05807_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07468__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07104__Y _02231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12765__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ clknet_leaf_85_clk _01281_ net1018 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10893__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13669_ clknet_leaf_86_clk _01228_ net1014 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08680__A2 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06210_ top.ru.state\[4\] top.busy_o top.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 _01427_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07190_ net808 net523 net463 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__o21a_1
XANTENNA_wire496_A _02779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12213__B1 _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07640__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09900_ _04881_ _04885_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09831_ net184 top.DUT.register\[1\]\[22\] net440 vssd1 vssd1 vccd1 vccd1 _00144_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout528 net529 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_4
Xfanout539 _03262_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06746__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10133__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ top.DUT.register\[13\]\[20\] net650 net550 top.DUT.register\[24\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a22o_1
X_09762_ top.pc\[16\] _04379_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__and2_1
XANTENNA__09207__B _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08111__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ _02120_ net489 net485 _02119_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a2bb2o_1
X_09693_ net344 _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08644_ _03334_ _03753_ _03754_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ _03687_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout443_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07459__A0 _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ top.DUT.register\[24\]\[4\] net551 net547 top.DUT.register\[5\]\[4\] _02643_
+ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11255__B2 top.a1.row2\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ top.DUT.register\[11\]\[6\] net642 net553 top.DUT.register\[7\]\[6\] _02583_
+ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a221o_1
XANTENNA__12435__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout708_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ _01496_ _01497_ net790 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_98_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12204__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _02508_ _02510_ _02512_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_98_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10375__Y _04950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ top.pc\[3\] _02739_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06339_ top.pad.button_control.debounce_dly top.pad.button_control.debounce vssd1
+ vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__and2b_2
XANTENNA__10308__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09058_ _01692_ _01734_ _01776_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06985__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ top.DUT.register\[2\]\[31\] net661 net547 top.DUT.register\[5\]\[31\] _03128_
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold560 top.DUT.register\[15\]\[30\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 top.DUT.register\[26\]\[21\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11020_ net30 net841 net811 net2145 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__o22a_1
Xhold582 top.DUT.register\[20\]\[31\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 top.DUT.register\[25\]\[25\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09923__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09687__A1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ clknet_leaf_29_clk _00535_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07698__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ _05754_ _05787_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07162__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11853_ _05688_ _05713_ _05694_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or3b_1
XANTENNA__09439__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10804_ net1533 net151 net353 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__mux2_1
X_11784_ _05624_ _05647_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11246__B2 top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ clknet_leaf_5_clk _01087_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ net156 net1769 net383 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08662__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07870__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ net2131 net175 net450 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
X_13454_ clknet_leaf_115_clk _01018_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12405_ clknet_leaf_90_clk _00041_ net998 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10218__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13385_ clknet_leaf_11_clk _00949_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10597_ net211 net1572 net387 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
XANTENNA__08414__A2 _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07875__X _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12336_ top.pad.button_control.r_counter\[4\] top.pad.button_control.r_counter\[3\]
+ _06126_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__and3_1
XANTENNA__07622__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06976__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12978__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ net891 top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__and2b_1
X_12198_ top.a1.row2\[17\] net846 net814 _06002_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__a22o_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ net132 _04624_ _05061_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__and3_1
XANTENNA_max_cap506_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10888__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07689__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__inv_2
XANTENNA__07153__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire509_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06900__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ _02636_ net469 _03480_ net482 _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07311_ top.DUT.register\[15\]\[9\] _01655_ net632 top.DUT.register\[19\]\[9\] _02437_
+ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a221o_1
X_08291_ _03413_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__nand2_2
XANTENNA__08653__A2 _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09850__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ top.DUT.register\[4\]\[14\] net769 net745 top.DUT.register\[31\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a22o_1
XANTENNA__07861__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06183__A_N top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ top.DUT.register\[28\]\[13\] net654 net553 top.DUT.register\[7\]\[13\] _02299_
+ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a221o_1
XANTENNA__10128__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07613__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11748__A top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout303 net309 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08122__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout325 _04957_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_6
XANTENNA__06719__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout336 net339 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_4
X_09814_ _04812_ _04813_ _04814_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__or3_1
Xfanout347 _04964_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_6
Xfanout358 net360 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1100_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _04958_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_6
X_09745_ _04740_ _04742_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__or3b_1
XANTENNA__10798__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ top.DUT.register\[10\]\[20\] net729 _02082_ _02083_ vssd1 vssd1 vccd1 vccd1
+ _02084_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout560_A _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ net259 net2294 net437 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__mux2_1
X_06888_ net513 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08627_ _03077_ _03736_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nand2_1
XANTENNA__13283__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A2 _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08558_ _02275_ _03664_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06864__X _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ _02634_ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__nand2_2
X_08489_ net317 _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10520_ net2193 net243 net363 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07852__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ net258 net1911 net369 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
XANTENNA__10038__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ clknet_leaf_49_clk _00734_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10382_ net151 net1998 net327 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
XANTENNA__06958__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ top.a1.dataIn\[3\] _05959_ _05960_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13404__RESET_B net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12052_ _05918_ _05920_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__o21a_1
Xhold390 top.DUT.register\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13646__Q net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ net1244 _05017_ net535 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__mux2_1
XANTENNA__08580__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 _01428_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08580__B2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout881 top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout892 top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_2
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06591__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__Y _01885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10501__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12954_ clknet_leaf_18_clk _00518_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06487__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 top.DUT.register\[19\]\[3\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12885_ clknet_leaf_5_clk _00449_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _05658_ _05677_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11767_ _05614_ _05635_ _05636_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a21oi_2
X_13506_ clknet_leaf_43_clk _01070_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10718_ net221 net1322 net383 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ _05540_ _05551_ _05559_ _05546_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13437_ clknet_leaf_104_clk _01001_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10649_ net1986 net244 net452 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08399__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13368_ clknet_leaf_16_clk _00932_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06950__A _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06949__A2 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net1392 _06118_ _06119_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_184_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13299_ clknet_leaf_3_clk _00863_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08213__Y _03339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12460__Q top.a1.instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09202__A_N _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ top.DUT.register\[5\]\[18\] net546 net598 top.DUT.register\[27\]\[18\] _02975_
+ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_166_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08020__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07374__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ top.DUT.register\[28\]\[24\] net653 net641 top.DUT.register\[11\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a22o_1
X_07791_ top.DUT.register\[10\]\[19\] net730 net718 top.DUT.register\[2\]\[19\] _02917_
+ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a221o_1
XANTENNA__06582__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09530_ top.pc\[27\] top.pc\[28\] _04532_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__and3_1
X_06742_ top.DUT.register\[17\]\[25\] net726 net673 top.DUT.register\[16\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
XANTENNA__10411__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _04488_ _04490_ _04487_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06673_ top.DUT.register\[15\]\[27\] _01655_ net631 top.DUT.register\[19\]\[27\]
+ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a221o_1
X_08412_ net285 _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09392_ _04434_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_195_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08343_ _02888_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout141_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _03394_ _03397_ net308 vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XANTENNA__09220__B _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ _02343_ _02345_ _02347_ _02351_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout406_A _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07156_ top.DUT.register\[6\]\[13\] net765 net749 top.DUT.register\[20\]\[13\] _02280_
+ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07087_ top.DUT.register\[20\]\[10\] net577 net623 top.DUT.register\[25\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a22o_1
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_4
XANTENNA_fanout775_A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08011__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout144 _04908_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_2
Xfanout155 _04900_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_1
Xfanout166 _04868_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
Xfanout177 net178 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_2
Xfanout188 _04820_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_1
XANTENNA_fanout942_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout199 net202 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ top.DUT.register\[26\]\[31\] net761 net672 top.DUT.register\[16\]\[31\] _03109_
+ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a221o_1
XANTENNA__06573__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ net207 net1906 net438 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XANTENNA__08314__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08314__B2 _03437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09659_ _02192_ _02193_ _02197_ _02203_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ clknet_leaf_14_clk _00234_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09411__A top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ _05474_ _05479_ _05483_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13029__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08617__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07825__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_1
Xwire512 _02099_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_2
Xwire523 _02316_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10503_ net184 net2320 net368 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11483_ _05338_ _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13222_ clknet_leaf_25_clk _00786_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10434_ net205 net1670 net325 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__mux2_1
XANTENNA__08461__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08314__X _03438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10365_ net1534 net157 net394 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ clknet_leaf_27_clk _00717_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08033__Y _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12104_ _05958_ _05969_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__xnor2_1
X_13084_ clknet_leaf_56_clk _00648_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10296_ net1546 net161 net401 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12035_ _05848_ _05904_ _05879_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08002__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__D _03875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08553__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__B1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__B2 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12538__RESET_B net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10231__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07106__A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ clknet_leaf_4_clk _00501_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09024__C _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12868_ clknet_leaf_39_clk _00432_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_199_Right_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ _05685_ _05686_ _05681_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09266__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ clknet_leaf_114_clk _00363_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07816__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07010_ top.DUT.register\[8\]\[11\] net742 net670 top.DUT.register\[5\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08224__X _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10406__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07595__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ net510 net591 net1206 net868 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ top.DUT.register\[6\]\[16\] net764 net708 top.DUT.register\[9\]\[16\] _03038_
+ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a221o_1
X_08892_ net522 _03985_ _03989_ net478 _03988_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__a221o_1
XANTENNA__07347__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12696__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08544__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06371__A_N top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _02961_ _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__nor2_8
XANTENNA__08400__A _03520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10351__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout189_A _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10141__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _02403_ _02900_ _02898_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_104_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09930__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07016__A _02142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09513_ top.pc\[27\] _04543_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_88_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06725_ top.DUT.register\[23\]\[26\] net562 net783 top.DUT.register\[31\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout356_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _04483_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__or2_1
X_06656_ top.DUT.register\[2\]\[27\] net719 net692 top.DUT.register\[21\]\[27\] _01780_
+ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ top.pc\[18\] _04394_ _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09257__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06587_ top.DUT.register\[19\]\[29\] net633 net787 top.DUT.register\[3\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08326_ _02685_ _02885_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07807__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08257_ _02783_ net468 _03380_ net476 _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__o221a_1
XFILLER_0_201_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08480__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07208_ top.DUT.register\[12\]\[15\] net580 net678 top.DUT.register\[13\]\[15\] _02334_
+ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a221o_1
X_08188_ _02682_ net289 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08134__X _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_A top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07139_ top.DUT.register\[21\]\[12\] net573 net656 top.DUT.register\[1\]\[12\] _02265_
+ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10316__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ net216 top.DUT.register\[8\]\[17\] net413 vssd1 vssd1 vccd1 vccd1 _00363_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ net229 net1596 net418 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__mux2_1
XANTENNA__07338__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09406__A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ net72 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ clknet_leaf_66_clk _01314_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10983_ top.a1.halfData\[3\] net798 net844 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ clknet_leaf_49_clk _00286_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ clknet_leaf_23_clk _00217_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__Y _03155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _05470_ _05471_ _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12584_ clknet_leaf_34_clk _00148_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11535_ _05403_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09750__A1_N net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__X _03171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11466_ _01391_ net267 _05297_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__a21o_1
X_13205_ clknet_leaf_6_clk _00769_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10417_ net260 net1779 net323 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__mux2_1
X_11397_ _05238_ _05256_ _05242_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10226__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07577__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ clknet_leaf_0_clk _00700_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10348_ net1739 net219 net394 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__mux2_1
XANTENNA__06785__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10279_ net1393 net224 net402 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__mux2_1
X_13067_ clknet_leaf_31_clk _00631_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07329__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09723__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ _05851_ _05879_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__o21a_1
X_13842__1111 vssd1 vssd1 vccd1 vccd1 _13842__1111/HI net1111 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_179_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10896__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06510_ top.a1.instruction\[20\] top.a1.instruction\[21\] net801 vssd1 vssd1 vccd1
+ vccd1 _01637_ sky130_fd_sc_hd__and3b_2
XFILLER_0_76_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07490_ top.DUT.register\[17\]\[5\] net643 net564 top.DUT.register\[4\]\[5\] _02616_
+ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06441_ net835 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09239__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09160_ _02608_ _02612_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__nor2_1
X_06372_ top.a1.instruction\[15\] top.a1.instruction\[16\] net810 vssd1 vssd1 vccd1
+ vccd1 _01499_ sky130_fd_sc_hd__and3b_2
XFILLER_0_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08111_ net318 net312 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09091_ _02205_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__nand2_1
XANTENNA__07777__Y _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13494__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09718__A1_N net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08042_ net296 net467 vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold901 top.DUT.register\[16\]\[17\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold912 top.DUT.register\[21\]\[10\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 top.DUT.register\[19\]\[9\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold934 top.DUT.register\[10\]\[29\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10136__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08974__A1_N net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 top.DUT.register\[24\]\[30\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07568__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 top.DUT.register\[8\]\[12\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 net43 vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 top.DUT.register\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold989 top.DUT.register\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net1799 net140 net432 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ top.pad.button_control.r_counter\[1\] top.pad.button_control.r_counter\[4\]
+ top.pad.button_control.r_counter\[3\] _04032_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_95_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1013_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11116__A3 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09714__B1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _03938_ _03955_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__o21a_1
X_07826_ top.DUT.register\[25\]\[18\] net774 net766 top.DUT.register\[6\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07757_ net298 net495 _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout640_A _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06708_ top.DUT.register\[17\]\[26\] net724 net677 top.DUT.register\[18\]\[26\] _01834_
+ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a221o_1
X_07688_ top.DUT.register\[2\]\[0\] net716 net681 top.DUT.register\[7\]\[0\] _02814_
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a221o_1
X_09427_ top.pc\[21\] _04434_ top.pc\[22\] vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a21oi_1
X_06639_ top.DUT.register\[23\]\[28\] net562 net618 top.DUT.register\[30\]\[28\] _01756_
+ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06700__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09358_ _04388_ _04391_ _04389_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_152_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ net320 _03432_ _03402_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_23_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08453__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09289_ _04337_ _04338_ _04339_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__o21ai_1
X_11320_ top.a1.dataIn\[22\] top.a1.dataIn\[21\] _05187_ top.a1.dataIn\[23\] vssd1
+ vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ top.a1.row1\[9\] _05108_ _05118_ top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1
+ _05130_ sky130_fd_sc_hd__a22o_1
XANTENNA__10046__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__A0 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__A0 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__B2 _03184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net264 net2230 net407 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
X_11182_ net1352 net533 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nand2b_1
X_10133_ net148 top.DUT.register\[8\]\[0\] net413 vssd1 vssd1 vccd1 vccd1 _00346_
+ sky130_fd_sc_hd__mux2_1
X_10064_ net464 _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__nand2_8
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_202_Right_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09181__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13367__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_67_clk _01364_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ clknet_leaf_91_clk _01297_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[43\]
+ sky130_fd_sc_hd__dfrtp_4
X_10966_ _01385_ net800 vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nand2_1
X_12705_ clknet_leaf_25_clk _00269_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13685_ clknet_leaf_95_clk _00016_ net990 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10897_ net2060 net160 net345 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12636_ clknet_leaf_17_clk _00200_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ clknet_leaf_106_clk _00131_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07798__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11518_ _05381_ _05387_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12498_ clknet_leaf_75_clk _00065_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold208 top.a1.data\[7\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold219 top.DUT.register\[28\]\[15\] vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13119_ clknet_leaf_114_clk _00683_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ _02102_ _02104_ _02115_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__nor4_2
X_08660_ net315 net480 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__nor2_2
XANTENNA__07183__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ _02207_ _02687_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08591_ _03507_ _03703_ net310 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_85_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06930__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07542_ top.DUT.register\[4\]\[4\] net768 net761 top.DUT.register\[26\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ top.DUT.register\[12\]\[5\] net580 net689 top.DUT.register\[3\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a22o_1
XANTENNA__13341__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08683__B1 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__Y _03989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ net137 _04256_ _04267_ net909 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__o211ai_1
X_06424_ top.DUT.register\[12\]\[30\] net581 net732 top.DUT.register\[19\]\[30\] _01550_
+ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__a221o_1
XANTENNA__12884__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06355_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__or4_1
X_09143_ _04201_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout221_A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout319_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07300__Y _02427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09074_ _01778_ _02123_ _02636_ _02685_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__or4bb_1
X_06286_ net1362 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[30\] sky130_fd_sc_hd__and2_1
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06997__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ _03150_ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__nor2_2
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold720 top.DUT.register\[31\]\[30\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold731 top.DUT.register\[15\]\[7\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold742 top.DUT.register\[23\]\[8\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08738__B2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 top.DUT.register\[4\]\[14\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold764 top.DUT.register\[1\]\[30\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold775 top.DUT.register\[14\]\[0\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06749__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 top.DUT.register\[23\]\[25\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap494 _02875_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_2
Xhold797 top.DUT.register\[1\]\[29\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ net1475 net195 net432 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
X_08927_ net318 _03726_ _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08858_ net2141 net840 net815 _03957_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_179_Left_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07174__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07713__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ top.DUT.register\[4\]\[19\] net566 net558 top.DUT.register\[6\]\[19\] _02935_
+ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__a221o_1
XANTENNA__06921__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ _01952_ _03177_ net485 _01950_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__a22o_1
XANTENNA__06586__Y _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ net1447 net227 net354 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11273__A2 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ net208 net1652 net375 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__C1 _04867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13470_ clknet_leaf_14_clk _01034_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ net240 net1993 net378 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10836__Y _04963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ clknet_leaf_94_clk top.ru.next_FetchedData\[5\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12352_ top.pad.button_control.r_counter\[9\] _06137_ top.pad.button_control.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08977__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__Q top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11303_ top.a1.row1\[15\] _05096_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12283_ _01445_ _06071_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11234_ _05092_ _05101_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13856__1121 vssd1 vssd1 vccd1 vccd1 _13856__1121/HI net1121 sky130_fd_sc_hd__conb_1
XANTENNA__10504__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ net1398 net532 net525 _05070_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ net1485 net212 net460 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
X_11096_ net914 net1294 net854 _05034_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ net228 net1640 net422 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__mux2_1
XANTENNA__07165__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06777__X _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 _01185_ vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold91 top.a1.data\[11\] vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06912__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13806_ clknet_leaf_64_clk _01349_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11998_ _05839_ _05865_ _05860_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__or3b_1
XFILLER_0_85_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ clknet_leaf_74_clk _01280_ net1018 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10949_ _01378_ _01418_ _01421_ _01410_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_158_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08665__B1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13668_ clknet_leaf_88_clk _01227_ net1007 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ clknet_leaf_29_clk _00183_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07768__B _02492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13599_ clknet_leaf_95_clk _01158_ net988 vssd1 vssd1 vccd1 vccd1 top.ramload\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06979__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10527__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09830_ _03864_ net340 net337 _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__o211a_4
Xfanout529 _01614_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_169_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07943__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ top.pc\[15\] _04362_ _04762_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_206_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ top.DUT.register\[19\]\[20\] net633 net787 top.DUT.register\[3\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a22o_1
X_08712_ _03817_ _03818_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__and2_1
X_09692_ top.a1.dataIn\[6\] _01492_ net803 top.pc\[6\] _04708_ vssd1 vssd1 vccd1 vccd1
+ _04709_ sky130_fd_sc_hd__a221o_1
XANTENNA__07156__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _03259_ _03741_ _03742_ net319 _03743_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__o221a_1
XANTENNA__06903__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08574_ net471 _03671_ _03673_ net475 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_25_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07459__A1 _02585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ top.DUT.register\[21\]\[4\] net575 net554 top.DUT.register\[7\]\[4\] _02651_
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_61_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ top.DUT.register\[2\]\[6\] net661 net570 top.DUT.register\[8\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06407_ top.DUT.register\[27\]\[30\] net776 net705 top.DUT.register\[15\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06682__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout603_A _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12204__B2 top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ top.DUT.register\[14\]\[7\] net721 net712 top.DUT.register\[30\]\[7\] _02513_
+ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_98_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ top.pc\[1\] _02788_ _04048_ _04047_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__a31o_1
XANTENNA__08959__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06338_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__and2_1
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06269_ net1320 net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[13\] sky130_fd_sc_hd__and2_1
X_09057_ _02781_ _03413_ _03523_ _03707_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08008_ top.DUT.register\[20\]\[31\] net578 net637 top.DUT.register\[16\]\[31\] _03134_
+ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a221o_1
Xhold550 top.DUT.register\[16\]\[25\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 top.DUT.register\[8\]\[24\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold572 top.DUT.register\[30\]\[30\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 top.DUT.register\[5\]\[20\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10324__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 top.DUT.register\[18\]\[30\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07934__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ net142 net2313 net435 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__mux2_1
X_12970_ clknet_leaf_34_clk _00534_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07147__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _05787_ _05789_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nor2_4
XFILLER_0_99_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11852_ _05679_ _05689_ net130 _05692_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10803_ net464 _04938_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_49_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08647__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _05641_ _05646_ _05649_ _05650_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__a211o_1
XFILLER_0_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13522_ clknet_leaf_50_clk _01086_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ net160 net1830 net381 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06673__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13453_ clknet_leaf_33_clk _01017_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10665_ net1335 net186 net452 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
X_12404_ clknet_leaf_82_clk _00040_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13384_ clknet_leaf_33_clk _00948_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ net217 net1927 net385 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12335_ _06128_ _06129_ net795 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and3b_1
XANTENNA__06425__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12266_ net2134 _06086_ net1107 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08052__X _03179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09375__A1 top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ net883 net885 vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or2_2
XFILLER_0_208_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10234__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
X_12197_ net2302 net846 net814 _06018_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__a22o_1
XANTENNA__07386__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__07925__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XANTENNA_output65_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ _04156_ _05060_ net897 _01618_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_182_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ net96 net862 net826 net1309 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07138__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13085__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07310_ top.DUT.register\[3\]\[9\] net786 net782 top.DUT.register\[31\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a22o_1
X_08290_ net312 _02731_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07310__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ top.DUT.register\[11\]\[14\] net757 net695 top.DUT.register\[21\]\[14\] _02367_
+ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a221o_1
XANTENNA__10409__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06664__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12198__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07172_ top.DUT.register\[14\]\[13\] net613 net610 top.DUT.register\[12\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_200_Left_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09281__A_N _02298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08403__A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09366__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10144__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net306 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
Xfanout315 net318 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07377__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 _04957_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_4
X_09813_ _04813_ _04814_ _04812_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09933__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
XANTENNA__07916__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout348 _04964_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_4
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_4
XANTENNA_fanout386_A _04945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__nand2_1
X_06956_ top.DUT.register\[22\]\[20\] net753 net742 top.DUT.register\[8\]\[20\] _02081_
+ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a221o_1
XANTENNA__07129__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13752__Q top.a1.row2\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _03391_ net341 net338 _04695_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__o211a_2
X_06887_ _02001_ _02006_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _03077_ _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout720_A _01527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _03669_ _03670_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout818_A _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07508_ _02608_ _02633_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__or2_1
X_08488_ _03386_ _03604_ net310 vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08137__X _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855__1120 vssd1 vssd1 vccd1 vccd1 _13855__1120/HI net1120 sky130_fd_sc_hd__conb_1
XANTENNA__10987__A1 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ top.a1.instruction\[27\] net528 _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06655__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12189__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ net259 net2035 net369 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _04154_ _04170_ _04145_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
XANTENNA__06407__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _01601_ _04937_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_60_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12120_ _05977_ _05984_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__xor2_1
XANTENNA__09409__A top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10054__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _05897_ _05898_ _05900_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09128__B _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 top.DUT.register\[9\]\[30\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold391 top.DUT.register\[7\]\[29\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ top.a1.dataIn\[9\] net848 net843 _05016_ vssd1 vssd1 vccd1 vccd1 _05017_
+ sky130_fd_sc_hd__a22o_1
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_2
Xfanout871 net873 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_2
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout893 top.a1.state\[0\] vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_2
X_12953_ clknet_leaf_37_clk _00517_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13662__Q net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1080 top.DUT.register\[6\]\[3\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 top.ramload\[15\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11904_ _05770_ _05771_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__or3_1
X_12884_ clknet_leaf_60_clk _00448_ net1099 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07540__B1 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__A top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11835_ _05689_ _05694_ _05696_ _05699_ _05703_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06894__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_185_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _05565_ _05612_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ clknet_leaf_27_clk _01069_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ net225 net2049 net382 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XANTENNA__10229__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _05550_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13436_ clknet_leaf_56_clk _01000_ net1086 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09045__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ net2180 net248 net450 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13367_ clknet_leaf_107_clk _00931_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10579_ net148 net2350 net385 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
X_12318_ top.lcd.cnt_500hz\[14\] _06118_ net588 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_184_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13298_ clknet_leaf_50_clk _00862_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12249_ _06071_ _06077_ net1108 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__o21a_1
XANTENNA__09038__B _03989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08020__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10899__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08571__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ top.DUT.register\[13\]\[24\] net647 net569 top.DUT.register\[8\]\[24\] _01932_
+ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a221o_1
X_07790_ top.DUT.register\[27\]\[19\] net777 net702 top.DUT.register\[29\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06741_ top.DUT.register\[28\]\[25\] net585 net748 top.DUT.register\[20\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ net906 top.pc\[23\] _04500_ net896 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__o211a_1
X_06672_ top.DUT.register\[3\]\[27\] net785 net781 top.DUT.register\[31\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a22o_1
XANTENNA__07531__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08411_ _03403_ _03408_ net299 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06885__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09391_ top.pc\[20\] _04413_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09808__C1 _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08342_ _02636_ _02887_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10969__A1 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ net286 _03301_ _03302_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__a31o_1
XANTENNA__06637__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout134_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09928__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07224_ top.DUT.register\[23\]\[15\] net560 net545 top.DUT.register\[5\]\[15\] _02350_
+ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07155_ top.DUT.register\[2\]\[13\] net717 net680 top.DUT.register\[13\]\[13\] _02281_
+ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout301_A _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ top.DUT.register\[13\]\[10\] net648 net612 top.DUT.register\[14\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a22o_1
XANTENNA__13747__Q top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
XANTENNA_fanout670_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 _04908_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_1
Xfanout156 _04890_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout768_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout167 _04868_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_1
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10602__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 _04840_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
Xfanout189 _04820_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
X_07988_ top.DUT.register\[11\]\[31\] net757 net724 top.DUT.register\[17\]\[31\] _03108_
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a221o_1
XFILLER_0_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12818__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ _03667_ net341 net338 _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__o211a_1
X_06939_ top.DUT.register\[3\]\[21\] net787 net783 top.DUT.register\[31\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ net465 _04680_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__nand2_8
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07522__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09251__X _04304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ net480 _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_106_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06876__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _04620_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11620_ _05488_ _05489_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _05375_ net250 _05417_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__o22a_2
XANTENNA__10049__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire502 _02446_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ net187 net2339 net367 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11482_ _05300_ net267 _05350_ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ clknet_leaf_116_clk _00785_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10433_ net213 top.DUT.register\[16\]\[18\] net326 vssd1 vssd1 vccd1 vccd1 _00620_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11385__A1 top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13152_ clknet_leaf_49_clk _00716_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07053__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08250__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13625__RESET_B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ net1467 net163 net393 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12561__Q top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12103_ _05965_ _05967_ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__nand3b_1
X_13083_ clknet_leaf_59_clk _00647_ net1098 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06800__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10295_ net1719 net164 net403 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
X_12034_ top.a1.dataIn\[4\] _05877_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09750__B2 top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06498__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 net691 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ clknet_leaf_31_clk _00500_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07106__B _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09024__D _03949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12867_ clknet_leaf_50_clk _00431_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11818_ _05681_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ clknet_leaf_15_clk _00362_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06619__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ _05602_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__or2_1
XANTENNA__09018__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07292__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ clknet_leaf_30_clk _00983_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_133_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07776__B _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07044__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08960_ _02231_ net591 net1185 net867 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11128__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ top.DUT.register\[22\]\[16\] net752 net705 top.DUT.register\[15\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__a22o_1
XANTENNA__06516__A_N top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net314 _03677_ _03745_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08544__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__A1 top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07842_ _02964_ _02966_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__or3_2
XFILLER_0_166_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10422__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07773_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_142_Left_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09512_ net907 top.pc\[26\] _04549_ net896 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_88_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06724_ top.DUT.register\[1\]\[26\] net657 net606 top.DUT.register\[18\]\[26\] _01850_
+ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09443_ top.pc\[23\] _04468_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06858__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06655_ top.DUT.register\[13\]\[27\] net678 net667 top.DUT.register\[5\]\[27\] _01781_
+ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout251_A _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_A _04963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ top.pc\[18\] _04394_ _04404_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06586_ _01704_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__nor2_8
XFILLER_0_191_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08128__A _03164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08325_ net313 _03447_ _03442_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11064__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07283__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ _02782_ _03177_ net484 _02781_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_151_Left_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ top.DUT.register\[1\]\[15\] net685 net674 top.DUT.register\[18\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08187_ _02731_ net294 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07035__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ top.DUT.register\[2\]\[12\] net660 net623 top.DUT.register\[25\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07069_ _01489_ _01491_ _01584_ _02187_ _02195_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__o221a_1
XANTENNA__07991__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ net180 net1894 net417 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10332__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13770_ clknet_leaf_66_clk _01313_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10982_ top.a1.dataInTemp\[3\] net800 vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ clknet_leaf_110_clk _00285_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06849__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12600__RESET_B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ clknet_leaf_10_clk _00216_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11603_ _05412_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_154_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ clknet_leaf_7_clk _00147_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11534_ _05348_ _05400_ _05389_ _05341_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08471__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06781__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ _01391_ _05297_ net267 vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__nand3_1
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13204_ clknet_leaf_47_clk _00768_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08759__C1 _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07026__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ net265 net1671 net325 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11396_ _05238_ _05242_ _05256_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ clknet_leaf_20_clk _00699_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10347_ net1370 net225 net396 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ clknet_leaf_38_clk _00630_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ net1857 net234 net401 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__mux2_1
X_12017_ _05852_ net127 _05859_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10242__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__B1 _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__C1 _04026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09332__A _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__B1 _01444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12919_ clknet_leaf_77_clk _00483_ net1085 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08388__A2_N _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06440_ net905 net904 top.a1.instruction\[6\] _01566_ vssd1 vssd1 vccd1 vccd1 _01567_
+ sky130_fd_sc_hd__nand4b_4
XTAP_TAPCELL_ROW_192_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12466__Q top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ top.a1.instruction\[17\] top.a1.instruction\[18\] net810 vssd1 vssd1 vccd1
+ vccd1 _01498_ sky130_fd_sc_hd__and3b_2
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ net316 net310 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__nor2_2
XFILLER_0_161_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09090_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__inv_2
XANTENNA__07265__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__A _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08041_ net291 net467 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_211_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10417__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold902 top.DUT.register\[6\]\[2\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold913 top.DUT.register\[4\]\[26\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 top.DUT.register\[18\]\[14\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold935 top.DUT.register\[16\]\[14\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 top.DUT.register\[23\]\[17\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold957 top.DUT.register\[20\]\[23\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 top.DUT.register\[6\]\[27\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ net1337 net144 net430 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
Xhold979 top.DUT.register\[17\]\[26\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08943_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[8\]
+ top.pad.button_control.r_counter\[6\] top.pad.button_control.r_counter\[2\] vssd1
+ vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__or4_1
XFILLER_0_209_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout299_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09714__B2 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08874_ net474 _03960_ _03972_ net471 _03970_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__o221a_1
XANTENNA__08130__B _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ top.DUT.register\[22\]\[18\] net754 net718 top.DUT.register\[2\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__a22o_1
XANTENNA__11772__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _02783_ _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nand2_1
X_06707_ top.DUT.register\[31\]\[26\] net746 net694 top.DUT.register\[21\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a22o_1
X_07687_ top.DUT.register\[22\]\[0\] net751 net689 top.DUT.register\[3\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout633_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ top.pc\[21\] top.pc\[22\] _04434_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__and3_1
X_06638_ top.DUT.register\[16\]\[28\] net637 net609 top.DUT.register\[12\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09357_ net139 _04402_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06569_ top.DUT.register\[4\]\[29\] net768 net706 top.DUT.register\[15\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _03431_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07256__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ net138 _04327_ _04334_ _01588_ net911 vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__o221a_1
XANTENNA__08453__B2 _03571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08239_ net272 _03358_ _03363_ net268 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10327__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07008__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11250_ net884 _05103_ net880 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__and3b_1
X_10201_ net148 net2303 net405 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
XANTENNA__08756__A2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _01407_ net533 _04636_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ net464 _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__nand2_4
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08321__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10063_ _04916_ _04921_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__nor2_4
XANTENNA__10062__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__C1 _04009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13822_ clknet_leaf_65_clk _01363_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13753_ clknet_leaf_91_clk _01296_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10965_ top.edg2.flip2 _04974_ top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__nor3b_2
X_12704_ clknet_leaf_44_clk _00268_ net1078 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13684_ clknet_leaf_92_clk _00015_ net990 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07495__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10896_ net1531 net164 net348 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ clknet_leaf_52_clk _00199_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06782__Y _01909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12566_ clknet_leaf_121_clk _00130_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07247__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__A1_N _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _05385_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10237__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12497_ clknet_leaf_75_clk _00064_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold209 top.DUT.register\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11448_ _05268_ _05303_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_189_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _05220_ _05221_ _05225_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__and3_1
X_13118_ clknet_leaf_13_clk _00682_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13049_ clknet_leaf_37_clk _00613_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12522__RESET_B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ _02207_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08590_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__inv_2
XANTENNA__08377__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07541_ top.DUT.register\[27\]\[4\] net777 _01535_ top.DUT.register\[3\]\[4\] _02667_
+ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07486__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ _02592_ _02593_ _02597_ _02598_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__or4_2
XANTENNA__08683__A1 _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08683__B2 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09211_ net133 _04261_ _04266_ net819 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__o22a_1
X_06423_ top.DUT.register\[13\]\[30\] net678 net675 top.DUT.register\[18\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09142_ top.pc\[4\] _02691_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__and2_1
X_06354_ _01482_ _01484_ vssd1 vssd1 vccd1 vccd1 top.ru.next_read_i sky130_fd_sc_hd__nor2_1
XANTENNA__07238__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09073_ _02494_ _04131_ _04132_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__or4b_1
X_06285_ net1363 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[29\] sky130_fd_sc_hd__and2_1
XANTENNA__10147__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout214_A _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ _03127_ _03148_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold710 top.DUT.register\[19\]\[14\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 top.DUT.register\[12\]\[25\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 top.DUT.register\[18\]\[27\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold743 top.DUT.register\[17\]\[4\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 top.DUT.register\[8\]\[7\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 top.DUT.register\[8\]\[26\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold776 top.DUT.register\[21\]\[24\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 top.DUT.register\[25\]\[5\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 top.DUT.register\[24\]\[27\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ net1833 net199 net431 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout583_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ net270 _03874_ _04021_ net269 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09699__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_X net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08857_ net886 top.pc\[27\] net539 _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout750_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07808_ top.DUT.register\[21\]\[19\] net575 net665 top.DUT.register\[29\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a22o_1
XANTENNA__10610__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ net316 _03565_ _03750_ net272 _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a221o_1
XFILLER_0_197_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ top.DUT.register\[6\]\[1\] net765 net582 top.DUT.register\[12\]\[1\] _02865_
+ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ net221 net2013 net375 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07477__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ top.pc\[21\] _04434_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ net244 net1862 net379 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ clknet_leaf_96_clk top.ru.next_FetchedData\[4\] net992 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[4\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07229__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_12351_ net1367 _06137_ _06139_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13051__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__D net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10057__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ top.a1.row1\[111\] _05161_ _05174_ _05098_ vssd1 vssd1 vccd1 vccd1 _05175_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ net1167 _06096_ _06097_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09387__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ net884 _05109_ net882 vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07937__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07401__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ top.a1.dataInTemp\[4\] top.a1.data\[4\] net799 vssd1 vssd1 vccd1 vccd1 _05070_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ top.DUT.register\[7\]\[17\] net216 net459 vssd1 vssd1 vccd1 vccd1 _00331_
+ sky130_fd_sc_hd__mux2_1
X_11095_ net69 net858 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__and2_1
X_10046_ net179 net1873 net421 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold70 top.a1.row1\[11\] vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 top.ramstore\[26\] vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10520__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 top.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13805_ clknet_leaf_64_clk _01348_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11997_ _05839_ net128 vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_67_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10948_ net844 _04977_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__nor2_2
XANTENNA__07468__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13736_ clknet_leaf_85_clk _01279_ net1018 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06676__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ clknet_leaf_87_clk _01226_ net1008 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10879_ net1458 net234 net346 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12618_ clknet_leaf_34_clk _00182_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13598_ clknet_leaf_95_clk _01157_ net988 vssd1 vssd1 vccd1 vccd1 top.ramload\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12213__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06428__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12549_ clknet_leaf_71_clk _00113_ net1095 vssd1 vssd1 vccd1 vccd1 top.a1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout519 net521 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12703__RESET_B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06600__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ top.a1.dataIn\[16\] net333 _04765_ net335 vssd1 vssd1 vccd1 vccd1 _04767_
+ sky130_fd_sc_hd__a211o_1
X_06972_ _02089_ _02093_ _02098_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_206_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__A1_N net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ _02122_ _03816_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__nand2_1
X_09691_ net836 _04227_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__nor2_1
Xfanout1090 net1092 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
X_08642_ _02909_ _03077_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__xor2_1
XANTENNA__10430__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ net480 _03676_ _03678_ net520 _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout164_A _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ top.DUT.register\[12\]\[4\] net609 net605 top.DUT.register\[18\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07455_ top.DUT.register\[28\]\[6\] net654 net565 top.DUT.register\[4\]\[6\] _02581_
+ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13207__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A _04920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06406_ _01497_ net790 _01508_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__and3_4
XFILLER_0_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07386_ top.DUT.register\[11\]\[7\] net755 net739 top.DUT.register\[8\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ net133 vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__inv_2
XANTENNA__06419__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06337_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__and2b_1
XFILLER_0_60_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07092__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _01993_ _02035_ _03920_ _03958_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__and4bb_1
X_06268_ net1287 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[12\] sky130_fd_sc_hd__and2_1
XFILLER_0_102_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_A _04969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08007_ top.DUT.register\[1\]\[31\] net657 net617 top.DUT.register\[30\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a22o_1
Xhold540 top.DUT.register\[16\]\[28\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10605__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06199_ top.a1.halfData\[0\] _01413_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__nor2_1
Xhold551 top.DUT.register\[5\]\[5\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 top.DUT.register\[3\]\[7\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 top.DUT.register\[8\]\[15\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold584 top.DUT.register\[16\]\[10\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 top.DUT.register\[26\]\[24\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_5_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ net144 net1868 net434 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__mux2_1
XANTENNA__09553__A_N _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ net268 _03496_ _03878_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _04869_ _04870_ _04871_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11920_ _05776_ _05783_ _05788_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a21o_1
XANTENNA__10340__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12121__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08895__B2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ _05681_ net130 _05715_ _05716_ _05719_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_185_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10802_ net1422 net141 net447 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ _05649_ _05651_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08647__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__B2 _03757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ net167 net1883 net383 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__mux2_1
XANTENNA__06658__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13521_ clknet_leaf_12_clk _01085_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_9_clk _01016_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10664_ net1529 net187 net452 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07870__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08046__A _03164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12403_ clknet_leaf_83_clk _00039_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_7_clk _00947_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10595_ net227 net2122 net386 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ top.pad.button_control.r_counter\[3\] _06126_ vssd1 vssd1 vccd1 vccd1 _06129_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07885__A _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08333__X _03456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07622__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06830__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ top.lcd.cnt_20ms\[11\] _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__and2_1
XANTENNA__12724__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10515__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11216_ net883 net885 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12196_ net1345 net846 net813 _06028_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__a22o_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XANTENNA__08583__B1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_208_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
X_11147_ _02789_ _02830_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ net1281 net862 net826 top.ramstore\[29\] vssd1 vssd1 vccd1 vccd1 _01196_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08335__B1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _04679_ _04921_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__nor2_2
XANTENNA__10250__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07689__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06897__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ clknet_leaf_67_clk _00002_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08227__Y _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10996__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07240_ top.DUT.register\[25\]\[14\] net774 net749 top.DUT.register\[20\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a22o_1
XANTENNA__07861__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12474__Q top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12198__A1 top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07171_ _02291_ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nor2_4
XFILLER_0_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12955__RESET_B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08390__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08810__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10425__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08403__B _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08574__B1 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout327 _04956_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_8
X_09812_ top.pc\[21\] _04460_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__nor2_1
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_4
Xfanout349 _04963_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_6
XANTENNA__09118__A2 _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ top.DUT.register\[28\]\[20\] net587 net758 top.DUT.register\[11\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a22o_1
X_09743_ top.pc\[14\] _04349_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout379_A _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10160__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ top.a1.dataIn\[2\] net794 net343 _04694_ vssd1 vssd1 vccd1 vccd1 _04695_
+ sky130_fd_sc_hd__a211o_1
X_06886_ _02008_ _02010_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_107_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08625_ _03709_ _03735_ _02359_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a21o_1
XANTENNA__11881__B1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ _02320_ _02904_ _03643_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_120_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07507_ _02608_ _02633_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__nand2_1
X_08487_ _03505_ _03603_ net304 vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout713_A _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_X net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10987__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07438_ _02206_ _02517_ _02564_ _01616_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_102_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09039__D1 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07852__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07369_ _02493_ _02494_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__nand2_2
X_09108_ net534 _04153_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ _04948_ _04953_ _04954_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__and3_2
XFILLER_0_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09039_ net316 _03559_ _03741_ net491 _03257_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06812__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ _05893_ _05896_ _05909_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__or4_1
Xhold370 top.DUT.register\[14\]\[22\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 top.DUT.register\[19\]\[7\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11001_ top.a1.data\[5\] top.a1.dataInTemp\[9\] net797 vssd1 vssd1 vccd1 vccd1 _05016_
+ sky130_fd_sc_hd__mux2_1
Xhold392 top.DUT.register\[25\]\[14\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout850 _04630_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_2
Xfanout861 _01430_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_2
Xfanout883 top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_2
Xfanout894 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_2
XANTENNA__06591__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10070__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ clknet_leaf_13_clk _00516_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08868__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1070 top.DUT.register\[10\]\[1\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 top.DUT.register\[18\]\[8\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09712__X _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1092 top.DUT.register\[24\]\[21\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ _05720_ _05765_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__xnor2_2
X_12883_ clknet_leaf_1_clk _00447_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08983__B _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _05696_ _05703_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09160__A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13522__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ _05621_ _05624_ _05625_ _05634_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13504_ clknet_leaf_44_clk _01068_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ net231 net1910 net382 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11696_ _05540_ _05559_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__and2_2
XANTENNA__09045__A1 _03350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10647_ net1647 net254 net451 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
X_13435_ clknet_leaf_57_clk _00999_ net1110 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ clknet_leaf_119_clk _00930_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10578_ net141 net1742 net358 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
XANTENNA__10245__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ _06118_ net588 _06117_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__and3b_1
X_13297_ clknet_leaf_118_clk _00861_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_197_Left_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ _06064_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap511_A _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12179_ _06047_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nand2_1
XANTENNA__08020__A2 _03146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08571__A3 _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06582__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ top.DUT.register\[10\]\[25\] net728 net690 top.DUT.register\[3\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06671_ top.DUT.register\[13\]\[27\] net647 net596 top.DUT.register\[27\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__a22o_1
X_08410_ net269 _03528_ _03529_ net272 _03527_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__a32o_1
XFILLER_0_176_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ top.pc\[20\] _04413_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__and2_1
XANTENNA__06694__A _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08341_ net1315 net837 net816 _03463_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a22o_1
XANTENNA__11615__B1 top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ net286 _03306_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07223_ top.DUT.register\[15\]\[15\] net779 _02348_ _02349_ vssd1 vssd1 vccd1 vccd1
+ _02350_ sky130_fd_sc_hd__a211o_1
XANTENNA__09036__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07047__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07154_ top.DUT.register\[22\]\[13\] net753 net670 top.DUT.register\[5\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
XANTENNA__09587__A2 _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07598__B2 top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10155__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07085_ net529 _02186_ _02211_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_2_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1036_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08011__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout135 _04185_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
Xfanout157 _04890_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_1
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout168 _04858_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_2
Xfanout179 net182 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
X_07987_ top.DUT.register\[8\]\[31\] net741 net714 top.DUT.register\[30\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout663_A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ _02058_ _02060_ _02062_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__or4_1
X_09726_ _04733_ _04734_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__o21ai_1
X_06869_ top.DUT.register\[20\]\[22\] net750 net746 top.DUT.register\[31\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
X_09657_ _04678_ _04679_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout928_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ net314 _03719_ _03718_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a21bo_1
X_09588_ top.pc\[31\] _04605_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08539_ net283 net298 _03203_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_46_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11550_ _05375_ _05379_ _05380_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__and3_1
XANTENNA__11082__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07825__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire503 _02423_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XFILLER_0_135_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ net193 net2227 net368 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__mux2_1
Xwire514 _02014_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_2
XFILLER_0_181_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ net267 _05299_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13220_ clknet_leaf_40_clk _00784_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10432_ net218 net2061 net323 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__mux2_1
X_13151_ clknet_leaf_111_clk _00715_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10363_ net1650 net166 net394 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10065__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08043__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ _05956_ _05964_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__xnor2_1
X_13082_ clknet_leaf_15_clk _00646_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ net1881 net168 net402 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
X_12033_ _05880_ _05901_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08002__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07210__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13673__Q top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout680 _01548_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_8
Xfanout691 _01541_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_70_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ clknet_leaf_7_clk _00499_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12866_ clknet_leaf_49_clk _00430_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11817_ _05685_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_194_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09266__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12797_ clknet_leaf_104_clk _00361_ net969 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11748_ top.a1.dataIn\[9\] _05589_ _05600_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__and3_1
XANTENNA__07816__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12547__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09018__A1 _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11679_ _05514_ _05547_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13418_ clknet_leaf_36_clk _00982_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_180_Right_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13349_ clknet_leaf_119_clk _00913_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08888__B _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ top.DUT.register\[28\]\[16\] net585 net668 top.DUT.register\[5\]\[16\] _03036_
+ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a221o_1
XANTENNA__10703__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ _01734_ net485 _03986_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a211o_1
X_07841_ top.DUT.register\[17\]\[18\] net725 net691 top.DUT.register\[3\]\[18\] _02967_
+ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a221o_1
XANTENNA__07201__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__A2 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _02298_ _02317_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__nand2b_1
X_06723_ top.DUT.register\[14\]\[26\] net613 net609 top.DUT.register\[12\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
X_09511_ net136 _04534_ _04548_ net907 vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06307__A2 _01445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ top.pc\[23\] _04468_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06654_ top.DUT.register\[26\]\[27\] net759 _01520_ top.DUT.register\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a22o_1
XANTENNA__08409__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09373_ _04416_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__nand2_1
XANTENNA__09257__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06585_ _01705_ _01707_ _01709_ _01711_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__or4_2
XFILLER_0_148_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08324_ _03409_ _03445_ _03444_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__a21o_1
XANTENNA__09939__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__Y _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08255_ _02783_ _03379_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ top.DUT.register\[28\]\[15\] net584 _02328_ _02332_ vssd1 vssd1 vccd1 vccd1
+ _02333_ sky130_fd_sc_hd__a211o_1
XANTENNA__07459__S net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08186_ _03303_ _03311_ net308 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07137_ top.DUT.register\[20\]\[12\] net578 net617 top.DUT.register\[30\]\[12\] _02263_
+ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a221o_1
X_07068_ _01476_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout780_A _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06794__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09709_ net236 net1715 net437 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
X_10981_ net1984 _05002_ net535 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12720_ clknet_leaf_122_clk _00284_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_143_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12651_ clknet_leaf_30_clk _00215_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_0__f_clk_X clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11602_ _05441_ _05442_ top.a1.dataIn\[13\] _05409_ vssd1 vssd1 vccd1 vccd1 _05472_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07259__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ clknet_leaf_19_clk _00146_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11533_ _05346_ _05401_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11464_ top.a1.dataIn\[16\] _05332_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10415_ net150 net2316 net323 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__mux2_1
X_13203_ clknet_leaf_1_clk _00767_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11395_ _05261_ _05263_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13134_ clknet_leaf_111_clk _00698_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10346_ net1558 net234 net395 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06785__A2 _01520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ clknet_leaf_4_clk _00629_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10277_ net2267 net236 net401 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__mux2_1
XANTENNA__10523__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _05867_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output40_A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ clknet_leaf_121_clk _00482_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07498__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09239__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12849_ clknet_leaf_110_clk _00413_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06370_ top.a1.instruction\[15\] top.a1.instruction\[16\] net810 vssd1 vssd1 vccd1
+ vccd1 _01497_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_83_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08040_ _03107_ _03152_ _03162_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_211_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold903 top.DUT.register\[28\]\[17\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 top.DUT.register\[24\]\[11\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 top.DUT.register\[26\]\[30\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 top.DUT.register\[9\]\[26\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 top.pad.keyCode\[1\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold958 top.DUT.register\[1\]\[26\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13390__CLK clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold969 top.DUT.register\[8\]\[14\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ net1473 net152 net431 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_11__f_clk_X clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10433__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ top.pad.button_control.r_counter\[16\] top.pad.button_control.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08480__A2_N net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ _03103_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout194_A _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07824_ _02949_ _02950_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__nor2_2
XANTENNA__09082__X _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ net288 _02875_ _02881_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout361_A _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06866__B _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout459_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ _01823_ _01825_ _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__or4_2
XANTENNA__07489__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ top.DUT.register\[28\]\[0\] net584 net667 top.DUT.register\[5\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a22o_1
XANTENNA__08139__A _01929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06637_ top.DUT.register\[21\]\[28\] net574 net649 top.DUT.register\[13\]\[28\] _01763_
+ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a221o_1
X_09425_ net906 top.pc\[21\] _04467_ net896 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06700__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09669__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09356_ top.pc\[18\] _04385_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__xnor2_1
X_06568_ top.DUT.register\[26\]\[29\] net761 net733 top.DUT.register\[19\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ net284 _03430_ _03407_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09287_ _04335_ _04336_ _04186_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_191_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06499_ net905 net904 _01476_ _01477_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10608__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08238_ _03361_ _03362_ net306 vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _03288_ _03294_ net299 vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10200_ net464 _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nand2_4
XFILLER_0_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ net1350 net532 net525 _05077_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _04685_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__nor2_2
XANTENNA__10343__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10062_ net141 net1593 net423 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13821_ clknet_leaf_63_clk _01362_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11276__A1 top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13752_ clknet_leaf_90_clk _01295_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_168_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ top.a1.row1\[63\] _04988_ _04979_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
XANTENNA__08049__A _03171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__X _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ clknet_leaf_115_clk _00267_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13683_ clknet_leaf_92_clk _00014_ net1000 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ net1648 net168 net346 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ clknet_leaf_18_clk _00198_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10518__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ clknet_leaf_6_clk _00129_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _05352_ _05373_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ clknet_4_13__leaf_clk _00063_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11447_ _05282_ _05310_ _05314_ _05315_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_111_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_189_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07404__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11378_ _05238_ _05243_ _05247_ _05229_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10329_ net1528 net167 net398 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__mux2_1
X_13117_ clknet_4_4__leaf_clk _00681_ net997 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10253__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12034__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07128__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ clknet_leaf_109_clk _00612_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07183__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06930__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07540_ top.DUT.register\[6\]\[4\] net765 _01514_ top.DUT.register\[16\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__B _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__Q top.a1.instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07471_ top.DUT.register\[22\]\[5\] net751 net743 top.DUT.register\[31\]\[5\] _02594_
+ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a221o_1
XFILLER_0_186_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08683__A2 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06422_ _01496_ _01499_ net792 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__and3_4
X_09210_ _04262_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07891__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12630__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ top.pc\[4\] _02691_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nor2_1
X_06353_ top.d_ready _01478_ _01481_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor3_1
XANTENNA__10428__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ _01735_ _01777_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__and3_1
XANTENNA__07643__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06284_ net1324 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[28\] sky130_fd_sc_hd__and2_1
XFILLER_0_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06997__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08023_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold700 top.DUT.register\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout207_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold711 top.DUT.register\[19\]\[29\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold722 top.DUT.register\[13\]\[31\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold733 top.DUT.register\[25\]\[31\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 top.DUT.register\[1\]\[31\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08422__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 top.DUT.register\[31\]\[31\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 top.DUT.register\[24\]\[10\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06749__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold777 top.DUT.register\[5\]\[30\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold788 top.DUT.register\[21\]\[27\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold799 top.DUT.register\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ net1402 net210 net432 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net307 _03947_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09699__A1 _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08856_ _03938_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__xor2_1
XFILLER_0_207_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07174__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09253__A _02142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ top.DUT.register\[13\]\[19\] net649 net621 top.DUT.register\[26\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a22o_1
X_08787_ net300 _03889_ _03887_ net269 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout743_A _01518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__C_N _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ top.DUT.register\[11\]\[1\] net757 net730 top.DUT.register\[10\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout910_A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07669_ top.DUT.register\[20\]\[0\] net576 net603 top.DUT.register\[18\]\[0\] _02795_
+ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09408_ net906 top.pc\[20\] _04437_ _04451_ net896 vssd1 vssd1 vccd1 vccd1 _00101_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07882__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12207__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ net249 net1714 net377 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ top.pc\[17\] _04370_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10338__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ top.pad.button_control.r_counter\[9\] _06137_ net796 vssd1 vssd1 vccd1 vccd1
+ _06139_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07634__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11301_ top.a1.row2\[15\] _05162_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or2_1
X_12281_ net1167 _06096_ net1107 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08603__Y _03715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ net880 _05096_ _05101_ net892 vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__and4b_2
XANTENNA__06404__X _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10073__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ net1339 net532 net525 _05069_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ net1435 net230 net461 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
X_11094_ net915 net1330 net854 _05033_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a31o_1
X_10045_ net197 net1849 net423 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__mux2_1
XANTENNA__10801__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08362__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 top.a1.dataInTemp\[11\] vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 top.pad.button_control.r_counter\[1\] vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 _01193_ vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 top.DUT.register\[25\]\[0\] vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06912__A2 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13804_ clknet_leaf_65_clk _01347_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11996_ _05825_ _05845_ _05839_ _05837_ _05836_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_58_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12653__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13735_ clknet_leaf_74_clk _01278_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10947_ _04977_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09862__A1 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__A2_N net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07873__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13666_ clknet_leaf_87_clk _01225_ net1008 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
X_10878_ net1539 net237 net345 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ clknet_leaf_3_clk _00181_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10248__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ clknet_leaf_98_clk _01156_ net984 vssd1 vssd1 vccd1 vccd1 top.ramload\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07625__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ clknet_leaf_79_clk _00112_ net1004 vssd1 vssd1 vccd1 vccd1 top.pc\[31\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__13179__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06979__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[31\] net997 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[31\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_2 _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09917__A2 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09057__B _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _02094_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_206_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _02122_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__or2_1
XANTENNA__10711__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ net247 net1978 net437 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__mux2_1
Xfanout1080 net1082 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07156__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ net273 _03750_ _03751_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__o21ai_4
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_2
XFILLER_0_174_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06903__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ _02320_ _03338_ _03685_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09801__A top.pc\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ top.DUT.register\[11\]\[4\] net641 net565 top.DUT.register\[4\]\[4\] _02649_
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout157_A _04890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10999__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07454_ top.DUT.register\[6\]\[6\] net559 net618 top.DUT.register\[30\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06405_ _01498_ net790 _01503_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__and3_1
XANTENNA__07321__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07385_ top.DUT.register\[12\]\[7\] net581 net728 top.DUT.register\[10\]\[7\] _02511_
+ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a221o_1
XANTENNA__10158__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout324_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06336_ top.pad.count\[1\] top.pad.count\[0\] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__and2b_1
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07616__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _01614_ _04175_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__nor2_1
XANTENNA__09947__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08813__C1 _03912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13531__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ _03735_ _03778_ _03815_ _03849_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__and4_1
X_06267_ net1252 net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[11\] sky130_fd_sc_hd__and2_1
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09369__B1 top.pc\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08006_ top.DUT.register\[6\]\[31\] net558 net609 top.DUT.register\[12\]\[31\] _03132_
+ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold530 top.DUT.register\[21\]\[19\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
X_06198_ _01419_ _01423_ _01422_ _01420_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[0\]
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_38_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout693_A _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 top.DUT.register\[27\]\[24\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 top.DUT.register\[19\]\[26\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold563 top.DUT.register\[14\]\[30\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 top.DUT.register\[20\]\[18\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 top.DUT.register\[24\]\[23\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 top.DUT.register\[17\]\[16\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ net152 net2344 net436 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ net522 _04004_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__nand2_1
XANTENNA__10621__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _04881_ _04882_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__nand2_1
XANTENNA__12484__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ net539 _03938_ _03939_ top.pc\[26\] net886 vssd1 vssd1 vccd1 vccd1 _03940_
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ _05681_ net130 _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__o21ai_2
X_10801_ net2041 net146 net446 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11781_ _05641_ _05646_ _05650_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a21o_1
XANTENNA__09844__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ clknet_leaf_0_clk _01084_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07855__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ net168 net1753 net382 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13451_ clknet_leaf_29_clk _01015_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10663_ net1598 net191 net452 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10068__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12402_ clknet_leaf_82_clk _00038_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ net181 net1474 net385 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
X_13382_ clknet_leaf_19_clk _00946_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12333_ top.pad.button_control.r_counter\[3\] _06126_ vssd1 vssd1 vccd1 vccd1 _06128_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07885__B _03011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_12264_ _06086_ net1107 _06085_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_186_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11215_ net891 net880 vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nor2_1
X_12195_ _06037_ _04976_ net846 net1291 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__a2bb2o_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__07386__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XANTENNA__09780__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__clkbuf_4
X_11146_ net132 _04624_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__clkbuf_4
XANTENNA__06594__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11077_ net93 net863 net827 net1198 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__a22o_1
XANTENNA__10531__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ net141 net1441 net426 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_201_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ top.a1.dataIn\[4\] _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nor2_1
XANTENNA__07846__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ clknet_leaf_67_clk _00001_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07310__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13649_ clknet_leaf_84_clk _01208_ net1017 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12198__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07170_ _02284_ _02285_ _02294_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__or4_4
XFILLER_0_171_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10706__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08810__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 net309 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07377__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
X_09811_ top.pc\[21\] _04460_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__and2_1
XANTENNA__08574__B2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout328 _04956_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
Xfanout339 _04688_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10441__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ top.pc\[14\] _04349_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__nand2_1
X_06954_ top.DUT.register\[19\]\[20\] net733 net699 top.DUT.register\[23\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a22o_1
XANTENNA__07129__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09673_ _01568_ net803 net895 vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__mux2_1
X_06885_ top.DUT.register\[29\]\[22\] net703 net672 top.DUT.register\[16\]\[22\] _02011_
+ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout274_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ _02360_ _02400_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08555_ _02904_ _03643_ _02320_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout441_A _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout539_A _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07506_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08486_ _03561_ _03602_ net277 vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_194_Right_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08147__A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__C1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07437_ _02207_ _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_A _01533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12189__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ _02494_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09107_ _04165_ _04168_ _04028_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06319_ _01331_ _01330_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__nor2_1
XANTENNA__08262__B1 _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_111_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07299_ _02206_ _02208_ _02425_ _01616_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__o211a_1
XANTENNA__10616__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09038_ _03375_ _03989_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08972__A1_N _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 top.DUT.register\[11\]\[26\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 top.DUT.register\[30\]\[26\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12665__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 top.lcd.currentState\[1\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10378__A_N net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold393 top.ramload\[4\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net1221 _05015_ net535 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__mux2_1
XANTENNA__06576__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _01493_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_4
Xfanout851 _04630_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_1
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_2
XANTENNA__10351__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 top.ru.next_iready vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_1
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_2
Xfanout895 top.pc\[2\] vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12951_ clknet_leaf_78_clk _00515_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1060 top.DUT.register\[9\]\[15\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 top.DUT.register\[15\]\[27\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ _05770_ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__nor2_1
Xhold1082 top.DUT.register\[4\]\[27\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 top.DUT.register\[10\]\[28\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ clknet_leaf_51_clk _00446_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07540__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ _05656_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09817__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07828__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09160__B _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ _05628_ _05633_ _05629_ _05632_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__or4b_1
XFILLER_0_68_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12575__Q top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13503_ clknet_leaf_114_clk _01067_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10715_ net236 net2086 net381 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11695_ _05561_ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ clknet_leaf_18_clk _00998_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ net1462 net256 net450 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__mux2_1
XANTENNA__09045__A2 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ clknet_leaf_6_clk _00929_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10526__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10577_ net145 net2331 net360 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\] _06114_ vssd1 vssd1 vccd1
+ vccd1 _06118_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ clknet_leaf_122_clk _00860_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08005__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ top.lcd.cnt_20ms\[3\] _06063_ top.lcd.cnt_20ms\[4\] vssd1 vssd1 vccd1 vccd1
+ _06076_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_75_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07359__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12178_ _06020_ _06045_ _06043_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_208_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10261__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ net56 net857 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09903__X _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06670_ _01790_ _01796_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__nor2_8
XANTENNA__13347__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07531__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08340_ net887 top.pc\[4\] net536 _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08271_ _03394_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__inv_2
XFILLER_0_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11105__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07222_ top.DUT.register\[31\]\[15\] net782 net619 top.DUT.register\[26\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__B net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07153_ top.DUT.register\[31\]\[13\] net745 net698 top.DUT.register\[23\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10436__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09441__C1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ _02208_ _02210_ _02207_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1029_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__A _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06558__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 net139 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 _04908_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
Xfanout158 _04890_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
XANTENNA__10171__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout169 _04858_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
X_07986_ top.DUT.register\[10\]\[31\] net730 net702 top.DUT.register\[29\]\[31\] _03112_
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ _04718_ _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__nor2_1
X_06937_ top.DUT.register\[23\]\[21\] net562 net558 top.DUT.register\[6\]\[21\] _02063_
+ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout656_A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ top.a1.instruction\[8\] _04675_ top.a1.instruction\[7\] vssd1 vssd1 vccd1
+ vccd1 _04679_ sky130_fd_sc_hd__nand3b_2
X_06868_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__inv_2
XANTENNA__07522__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ net284 net299 _03429_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or3_2
XFILLER_0_179_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09587_ top.pc\[30\] _04587_ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a21o_1
XANTENNA__06730__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ top.DUT.register\[11\]\[24\] net757 net695 top.DUT.register\[21\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _02276_ net488 vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ _02448_ net488 net486 _02449_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08483__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire504 _02357_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_2
X_10500_ net206 net1590 net367 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire515 _01948_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_2
X_11480_ _05257_ _05298_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10431_ net228 net2002 net324 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10346__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ clknet_leaf_13_clk _00714_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ net1433 net170 net396 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06797__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _05969_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13081_ clknet_leaf_34_clk _00645_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10293_ net1727 net173 net403 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12032_ _05901_ _05880_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06412__X _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 top.a1.row1\[123\] vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06549__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09155__B _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _01554_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_4
Xfanout681 net684 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_8
Xfanout692 _01540_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12934_ clknet_leaf_19_clk _00498_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08339__X _03462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ clknet_leaf_27_clk _00429_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06721__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11206__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ _05642_ _05682_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_194_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12796_ clknet_leaf_17_clk _00360_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_194_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _05592_ _05601_ _05615_ _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_166_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09018__A2 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11678_ _05514_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ clknet_leaf_4_clk _00981_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10256__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10629_ net213 top.DUT.register\[22\]\[18\] net392 vssd1 vssd1 vccd1 vccd1 _00812_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08777__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13348_ clknet_leaf_39_clk _00912_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06788__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ clknet_leaf_113_clk _00843_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_47_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11128__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07840_ top.DUT.register\[23\]\[18\] net699 net680 top.DUT.register\[13\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__a22o_1
XANTENNA_max_cap507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07771_ _02399_ _02380_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06960__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ net132 _04538_ _04539_ _04547_ net819 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__o32a_1
X_06722_ top.DUT.register\[21\]\[26\] net574 net601 top.DUT.register\[10\]\[26\] _01848_
+ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13375__RESET_B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09441_ net906 top.pc\[22\] _04482_ net896 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__o211a_1
X_06653_ top.DUT.register\[20\]\[27\] net747 net727 top.DUT.register\[10\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_56_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ top.pc\[19\] _04407_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06584_ top.DUT.register\[29\]\[29\] net702 net682 top.DUT.register\[7\]\[29\] _01710_
+ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a221o_1
X_08323_ _03444_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08254_ _02877_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08425__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07205_ top.DUT.register\[26\]\[15\] net759 net704 top.DUT.register\[15\]\[15\] _02327_
+ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a221o_1
X_08185_ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout404_A _04939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09955__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__X _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ top.DUT.register\[13\]\[12\] net649 net602 top.DUT.register\[10\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07067_ net904 _01481_ top.a1.instruction\[4\] vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07991__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09690__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ _03089_ _03094_ _01953_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _03571_ net341 net338 _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o211a_2
X_10980_ top.a1.dataIn\[2\] net849 _04999_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_74_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07504__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09639_ top.a1.halfData\[2\] _01472_ _04665_ net1103 vssd1 vssd1 vccd1 vccd1 _00118_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06703__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ clknet_leaf_34_clk _00214_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ top.a1.dataIn\[12\] _05444_ _05445_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__or3_1
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ clknet_leaf_120_clk _00145_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_176_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11532_ _05346_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10076__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13042__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ _05325_ _05329_ _05331_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08759__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13202_ clknet_leaf_51_clk _00766_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10414_ _04686_ _04955_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_59_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11394_ _05261_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__nor2_1
X_13133_ clknet_leaf_32_clk _00697_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10804__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ net1509 net238 net393 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ clknet_leaf_34_clk _00628_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ net1801 net239 net402 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ _05865_ net127 _05860_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__and3b_1
XANTENNA__09723__A3 _04318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08931__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__B2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06942__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07414__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12917_ clknet_leaf_6_clk _00481_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09892__C1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12848_ clknet_leaf_0_clk _00412_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ clknet_leaf_31_clk _00343_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold904 top.DUT.register\[25\]\[7\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold915 top.DUT.register\[17\]\[6\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold926 top.DUT.register\[25\]\[8\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 top.DUT.register\[28\]\[25\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold948 top.DUT.register\[29\]\[13\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ net1909 net156 net431 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__mux2_1
XANTENNA__10714__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold959 top.DUT.register\[21\]\[9\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09076__A _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _04032_ _04035_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__nor2_1
XANTENNA__11506__B1 top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08872_ _01778_ _03102_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_209_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07186__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07725__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ _02928_ _02948_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06933__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout187_A _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07754_ _02831_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06705_ top.DUT.register\[27\]\[26\] net777 net741 top.DUT.register\[8\]\[26\] _01829_
+ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07685_ top.DUT.register\[12\]\[0\] net580 net755 top.DUT.register\[11\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
XANTENNA__08686__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout354_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1096_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09424_ net136 _04452_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__o21ai_1
X_06636_ top.DUT.register\[29\]\[28\] net665 net622 top.DUT.register\[26\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09355_ net907 top.pc\[17\] _04401_ net896 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__o211a_1
XANTENNA__12376__S _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06567_ _01692_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__nor2_2
XFILLER_0_118_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ _03408_ _03429_ net299 vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09286_ _04335_ _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__and2_1
XANTENNA__08155__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06498_ net805 _01623_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__or2_2
XFILLER_0_191_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09650__A2 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ _03225_ _03232_ net287 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09685__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ _03292_ _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07119_ top.DUT.register\[9\]\[12\] net709 net676 top.DUT.register\[18\]\[12\] _02245_
+ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a221o_1
XANTENNA__10624__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ net289 _02875_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__nand2_1
X_10130_ top.a1.instruction\[9\] top.a1.instruction\[10\] _04675_ vssd1 vssd1 vccd1
+ vccd1 _04929_ sky130_fd_sc_hd__nand3b_4
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09166__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ net147 net1937 net422 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
XANTENNA__07177__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__B2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06924__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_63_clk _01361_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07505__Y _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ clknet_leaf_88_clk _01294_ net1005 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[40\]
+ sky130_fd_sc_hd__dfrtp_2
X_10963_ top.a1.halfData\[0\] _01415_ _01417_ top.a1.hexop\[3\] net849 vssd1 vssd1
+ vccd1 vccd1 _04988_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12702_ clknet_leaf_13_clk _00266_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13682_ clknet_leaf_94_clk _00013_ net993 vssd1 vssd1 vccd1 vccd1 top.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894_ net1898 net173 net347 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12633_ clknet_leaf_35_clk _00197_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12861__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12564_ clknet_leaf_60_clk _00128_ net1099 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08065__A _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07101__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11515_ _05361_ _05383_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12495_ clknet_leaf_45_clk _00062_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramstore\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _05314_ _05315_ _05312_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10534__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11200__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11377_ _05199_ _05245_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ clknet_leaf_56_clk _00680_ net1086 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ net1625 net169 net398 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13047_ clknet_leaf_105_clk _00611_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ net2016 net169 net455 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__mux2_1
XANTENNA__07168__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07415__Y _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08668__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__A2 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10475__A0 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ top.DUT.register\[1\]\[5\] net685 net678 top.DUT.register\[13\]\[5\] _02595_
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07340__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06421_ net790 _01503_ _01508_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12216__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10709__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _04187_ _04190_ _04189_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__a21o_1
X_06352_ _01483_ vssd1 vssd1 vccd1 vccd1 top.ru.next_write_i sky130_fd_sc_hd__inv_2
XFILLER_0_127_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06283_ net1325 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[27\] sky130_fd_sc_hd__and2_1
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11113__B net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09071_ _01693_ _01907_ _03076_ _03151_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__and4_1
XANTENNA__08840__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ net490 _03147_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold701 top.DUT.register\[7\]\[15\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 top.DUT.register\[22\]\[31\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 top.DUT.register\[25\]\[26\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold734 top.DUT.register\[6\]\[15\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10444__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold745 top.DUT.register\[22\]\[21\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08422__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold756 top.DUT.register\[15\]\[6\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 top.DUT.register\[21\]\[17\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 _03072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 top.DUT.register\[22\]\[13\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ net2346 net219 net431 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_139_Left_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_1
Xhold789 top.DUT.register\[5\]\[3\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09148__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ net281 _03980_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07159__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _01818_ net489 _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__o21a_2
XANTENNA_fanout471_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ top.DUT.register\[23\]\[19\] net563 net597 top.DUT.register\[27\]\[19\] _02932_
+ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a221o_1
XANTENNA__09253__B _04304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ _03856_ _03888_ net277 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07737_ top.DUT.register\[28\]\[1\] net586 net683 top.DUT.register\[7\]\[1\] _02863_
+ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout736_A _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07668_ top.DUT.register\[11\]\[0\] net639 net619 top.DUT.register\[26\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_148_Left_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07331__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09407_ _04186_ _04442_ _04448_ _04450_ _01386_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a221o_1
X_06619_ top.DUT.register\[12\]\[28\] net582 net676 top.DUT.register\[18\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a22o_1
XANTENNA__12207__A1 top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10619__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A top.a1.instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ top.DUT.register\[28\]\[3\] net584 net712 top.DUT.register\[30\]\[3\] _02725_
+ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11304__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ top.pc\[17\] _04370_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__and2_1
XANTENNA__09084__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08831__B1 _03878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _04319_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11300_ net1203 net824 _05173_ net1095 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__o211a_1
X_12280_ _06096_ net1107 _06095_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__and3b_1
XFILLER_0_160_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09387__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ _05097_ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__nor2_1
XANTENNA__10354__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ top.a1.data\[3\] net797 _05003_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__o21a_1
XANTENNA__13407__RESET_B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ net1861 net179 net459 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11093_ net68 net858 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__and2_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net200 net1638 net423 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
XANTENNA__08898__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 top.ramstore\[13\] vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A2 _03483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 top.a1.data\[8\] vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 _01354_ vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold83 top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 net95 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07570__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13803_ clknet_leaf_64_clk _01346_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11249__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11995_ _05861_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13734_ clknet_leaf_74_clk _01277_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10946_ _04974_ net814 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__or2_2
XFILLER_0_202_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06676__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13665_ clknet_leaf_86_clk _01224_ net1007 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
X_10877_ net1928 net239 net345 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__mux2_1
XANTENNA__10529__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ clknet_leaf_32_clk _00180_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13596_ clknet_leaf_95_clk _01155_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12547_ clknet_leaf_79_clk _00111_ net1013 vssd1 vssd1 vccd1 vccd1 top.pc\[30\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06428__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ clknet_leaf_95_clk top.ru.next_FetchedInstr\[30\] net991 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[30\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_3 top.ru.next_FetchedData\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11429_ _05257_ _05295_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__xor2_1
XANTENNA__10264__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07928__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08810__X _03912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06600__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06970_ top.DUT.register\[26\]\[20\] net762 net672 top.DUT.register\[16\]\[20\] _02090_
+ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_169_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08889__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1076 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_2
X_08640_ _03186_ _03542_ _03564_ net271 vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__o22a_1
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_175_Right_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1092 net1097 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XFILLER_0_174_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ net320 net522 _03683_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_46_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_178_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07522_ top.DUT.register\[6\]\[4\] net559 net614 top.DUT.register\[14\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08257__X _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07313__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10999__A1 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07453_ _02571_ _02573_ _02575_ _02579_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__or4_1
XANTENNA__06667__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06404_ _01499_ net792 _01508_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__and3_4
XFILLER_0_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07321__B _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ top.DUT.register\[31\]\[7\] net744 net680 top.DUT.register\[13\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09123_ net137 _04182_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_98_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06335_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__nor2_1
XANTENNA__06419__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1059_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _04078_ _04079_ _04085_ _04086_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06266_ net2111 net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[10\] sky130_fd_sc_hd__and2_1
XANTENNA__07092__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09369__A1 top.pc\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ top.DUT.register\[24\]\[31\] net550 net621 top.DUT.register\[26\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a22o_1
Xhold520 top.DUT.register\[9\]\[22\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10174__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06197_ top.a1.hexop\[2\] top.a1.hexop\[3\] top.a1.hexop\[4\] vssd1 vssd1 vccd1 vccd1
+ _01423_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_38_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold531 top.DUT.register\[10\]\[3\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold542 top.DUT.register\[29\]\[7\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11176__B2 _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 top.DUT.register\[12\]\[20\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 top.DUT.register\[13\]\[18\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 top.DUT.register\[29\]\[11\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold586 top.DUT.register\[9\]\[19\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 top.DUT.register\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ net156 net2150 net435 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
XANTENNA__06888__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ net322 _03704_ _03859_ net271 _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o221a_1
X_09887_ top.pc\[28\] _04578_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10687__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _03916_ _03937_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07552__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _03839_ _03872_ net282 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_169_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10800_ net1686 net154 net447 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__mux2_1
X_11780_ _05617_ _05639_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07304__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10731_ net172 net1997 net384 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
XANTENNA__06658__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10349__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ clknet_leaf_38_clk _01014_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10662_ net1692 net204 net451 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ clknet_leaf_82_clk _00037_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07607__B2 top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ clknet_leaf_119_clk _00945_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10593_ net195 top.DUT.register\[21\]\[14\] net388 vssd1 vssd1 vccd1 vccd1 _00776_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12332_ _06126_ _06127_ net795 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__and3b_1
XFILLER_0_106_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ top.lcd.cnt_20ms\[10\] top.lcd.cnt_20ms\[9\] _06082_ vssd1 vssd1 vccd1 vccd1
+ _06086_ sky130_fd_sc_hd__and3_1
XANTENNA__06830__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11214_ _05092_ _05093_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__and2b_1
X_12194_ net1327 net846 net813 _06045_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__a22o_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__08583__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__A1 _03776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_11145_ _01448_ _01468_ _01469_ _01449_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__o211a_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10812__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__07791__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ net1217 net856 net825 top.ramstore\[27\] vssd1 vssd1 vccd1 vccd1 _01194_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08335__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net145 net1875 net428 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07543__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06897__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_201_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ _05752_ _05846_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13717_ clknet_leaf_67_clk _00000_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10929_ net165 net1941 net443 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XANTENNA__10259__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13648_ clknet_leaf_87_clk _01207_ net1005 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13579_ clknet_leaf_95_clk _01138_ net990 vssd1 vssd1 vccd1 vccd1 top.ramload\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08540__X _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
X_09810_ _04803_ _04805_ _04804_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a21oi_1
Xfanout318 _02663_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10722__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08700__B net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ top.a1.dataIn\[14\] _04720_ _04749_ _04718_ vssd1 vssd1 vccd1 vccd1 _04750_
+ sky130_fd_sc_hd__a211o_1
X_06953_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__inv_2
XANTENNA__12222__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09523__A1 _01840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ net266 net1513 net439 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__mux2_1
X_06884_ top.DUT.register\[26\]\[22\] net761 net682 top.DUT.register\[7\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09812__A top.pc\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ net1786 net840 net815 _03734_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_19_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08554_ net1493 net840 net815 _03668_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a22o_1
XANTENNA__09287__B1 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07505_ net805 _02612_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__o21ai_4
X_08485_ _03246_ _03250_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__nand2_1
XANTENNA__10169__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout434_A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08147__B net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09958__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ top.a1.instruction\[18\] net524 _01621_ top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09039__B1 _03741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout601_A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07367_ net499 _02492_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__nand2_1
X_09106_ _04164_ net534 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__nand2b_1
X_06318_ net1106 _01451_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08262__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08163__A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07298_ _02207_ _02424_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ _03879_ _03950_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__nand2_1
X_06249_ net1497 net873 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[25\] sky130_fd_sc_hd__and2_1
XANTENNA__06812__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_211_Right_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold350 top.DUT.register\[28\]\[29\] vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout970_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 top.DUT.register\[7\]\[7\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 top.DUT.register\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 top.DUT.register\[24\]\[20\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10632__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 top.DUT.register\[20\]\[24\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout830 _05024_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_2
Xfanout841 _05023_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_2
Xfanout852 net855 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07507__A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ net219 net2009 net435 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__mux2_1
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_181_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 top.ru.next_iready vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_2
Xfanout885 top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_2
Xfanout896 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_4
X_12950_ clknet_leaf_121_clk _00514_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1050 top.DUT.register\[21\]\[7\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1061 top.DUT.register\[24\]\[22\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _05727_ _05768_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1072 top.DUT.register\[18\]\[25\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 top.DUT.register\[18\]\[23\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ clknet_leaf_118_clk _00445_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1094 top.DUT.register\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11832_ _05654_ _05700_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_64_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13149__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11763_ _05572_ _05604_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__xor2_2
XFILLER_0_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10079__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13502_ clknet_leaf_10_clk _01066_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10714_ net240 net2064 net382 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11694_ _05552_ _05558_ _05557_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13433_ clknet_leaf_37_clk _00997_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ net1783 net262 net450 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
XANTENNA__10807__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ clknet_leaf_46_clk _00928_ net1083 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10576_ net154 top.DUT.register\[20\]\[29\] net358 vssd1 vssd1 vccd1 vccd1 _00759_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12315_ top.lcd.cnt_500hz\[12\] _01439_ _06109_ top.lcd.cnt_500hz\[13\] vssd1 vssd1
+ vccd1 vccd1 _06117_ sky130_fd_sc_hd__a31o_1
X_13295_ clknet_leaf_19_clk _00859_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12246_ _06071_ _06075_ net1108 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10542__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _06019_ _06043_ _06045_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_166_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11128_ net918 net1166 net852 _05050_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11059_ net74 net860 net829 net1185 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a22o_1
XANTENNA__07516__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09808__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ net280 _03298_ _03299_ _03393_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07221_ top.DUT.register\[19\]\[15\] net632 net785 top.DUT.register\[3\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__a22o_1
XANTENNA__10717__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07047__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ _02236_ _02277_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07083_ _01387_ _01616_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13858__1149 vssd1 vssd1 vccd1 vccd1 net1149 _13858__1149/LO sky130_fd_sc_hd__conb_1
XANTENNA__10452__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
Xfanout159 _04890_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_1
X_07985_ top.DUT.register\[23\]\[31\] net699 net694 top.DUT.register\[21\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout384_A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ net835 _04312_ _04720_ top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 _04735_
+ sky130_fd_sc_hd__a2bb2o_1
X_06936_ top.DUT.register\[1\]\[21\] net658 net622 top.DUT.register\[26\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a22o_1
X_09655_ top.a1.instruction\[9\] top.a1.instruction\[10\] _04675_ vssd1 vssd1 vccd1
+ vccd1 _04678_ sky130_fd_sc_hd__o21a_2
X_06867_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__or2_2
XFILLER_0_179_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout551_A _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ net268 _03527_ _03531_ net272 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a22oi_2
XANTENNA_fanout649_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_09586_ top.pc\[30\] _04587_ _04611_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__o21a_1
X_06798_ top.DUT.register\[14\]\[24\] net723 net700 top.DUT.register\[29\]\[24\] _01924_
+ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08537_ net317 _03651_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08468_ _03295_ _03541_ _03576_ net319 _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__a221oi_2
XANTENNA__09680__A0 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11082__A3 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ top.DUT.register\[25\]\[6\] net773 net694 top.DUT.register\[21\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
Xwire505 _02273_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ net472 _03493_ _03513_ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10430_ net179 net1617 net323 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ net1387 net171 net395 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12100_ _05940_ _05968_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07994__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ clknet_leaf_108_clk _00644_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10292_ net2017 net175 net401 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XANTENNA__08621__A _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _05886_ _05888_ _05894_ _05899_ _05883_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__o41a_2
Xhold180 top.ramload\[0\] vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10362__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 top.ramstore\[5\] vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07210__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 _01638_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_2
Xfanout671 net673 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_8
Xfanout682 net683 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_8
Xfanout693 _01540_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__Y _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ clknet_leaf_120_clk _00497_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09171__B _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12864_ clknet_leaf_45_clk _00428_ net1082 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08068__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11058__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11815_ top.a1.dataIn\[6\] _05682_ _05683_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ clknet_leaf_57_clk _00359_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_194_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13674__RESET_B net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ top.a1.dataIn\[9\] _05528_ _05560_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09671__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10537__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _05512_ _05541_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11222__A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07029__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13416_ clknet_leaf_32_clk _00980_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10628_ net215 net2336 net389 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08226__B2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13347_ clknet_leaf_50_clk _00911_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09974__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10559_ net208 net2021 net358 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__mux2_1
XANTENNA__07985__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ clknet_leaf_13_clk _00842_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12229_ net1220 _05975_ net589 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_102_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10272__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07737__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07201__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07770_ _02339_ _02358_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__nand2b_1
X_06721_ top.DUT.register\[28\]\[26\] net653 net645 top.DUT.register\[17\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XANTENNA__09362__A _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09440_ net132 _04475_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08701__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06652_ top.DUT.register\[6\]\[27\] net763 net751 top.DUT.register\[22\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11049__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09371_ top.pc\[19\] _04407_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_111_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06583_ top.DUT.register\[14\]\[29\] net722 net709 top.DUT.register\[9\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08971__A1_N _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ net298 _03203_ net283 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ _02878_ _03170_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08425__B net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07204_ _02324_ _02325_ _02329_ _02330_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__or4_2
XFILLER_0_144_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08184_ _03306_ _03309_ net280 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07135_ top.DUT.register\[4\]\[12\] net566 net542 top.DUT.register\[22\]\[12\] _02261_
+ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07066_ _01495_ net524 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout599_A _01669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__A0 _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _03089_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06919_ top.DUT.register\[20\]\[21\] net750 net746 top.DUT.register\[31\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a22o_1
X_09707_ top.pc\[8\] net803 _04718_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a211o_1
X_07899_ top.DUT.register\[16\]\[17\] net635 net781 top.DUT.register\[31\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _04659_ _04663_ _04664_ _04654_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__or4b_1
XANTENNA__07504__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ top.pc\[29\] _04566_ top.pc\[30\] vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ _05409_ _05444_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ clknet_leaf_39_clk _00144_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07259__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11531_ _05372_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__and2_1
XANTENNA__10357__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11462_ _05325_ _05329_ _05331_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ clknet_leaf_110_clk _00765_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10413_ net140 net2014 net330 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__mux2_1
X_11393_ _05237_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_59_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13132_ clknet_leaf_8_clk _00696_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10344_ net1877 net242 net393 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__mux2_1
XANTENNA__07431__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09708__A1 _03571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10092__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ clknet_leaf_8_clk _00627_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10275_ net2198 net245 net404 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07719__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _05860_ _05861_ net127 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__and3_1
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10820__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 net492 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_4
XANTENNA__11217__A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ clknet_leaf_60_clk _00480_ net1102 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07414__B _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ clknet_leaf_22_clk _00411_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857__1148 vssd1 vssd1 vccd1 vccd1 net1148 _13857__1148/LO sky130_fd_sc_hd__conb_1
X_12778_ clknet_leaf_40_clk _00342_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11223__Y _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11729_ _05595_ _05597_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold905 top.DUT.register\[16\]\[8\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold916 top.DUT.register\[28\]\[30\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 top.DUT.register\[18\]\[11\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09357__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 top.DUT.register\[26\]\[18\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold949 top.DUT.register\[10\]\[6\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06630__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ top.pad.button_control.r_counter\[8\] _04034_ top.pad.button_control.r_counter\[10\]
+ top.pad.button_control.r_counter\[9\] vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__o211a_1
XANTENNA__09076__B _01865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08871_ _03654_ _03771_ _03963_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_209_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07822_ _02928_ _02948_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__and2_1
XFILLER_0_209_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10730__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__X _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _02879_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__inv_2
XANTENNA__12854__CLK clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ top.DUT.register\[22\]\[26\] net753 net679 top.DUT.register\[13\]\[26\] _01830_
+ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07489__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ net805 _02788_ _02809_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ net132 _04458_ _04464_ _04465_ net906 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o221a_1
XFILLER_0_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06635_ top.DUT.register\[11\]\[28\] net641 net558 top.DUT.register\[6\]\[28\] _01761_
+ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a221o_1
XANTENNA__06697__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09820__A top.pc\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09354_ net136 _04387_ _04400_ net906 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout1089_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06566_ _01560_ _01690_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06508__X _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ net282 _03347_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09285_ _04313_ _04314_ _04315_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10177__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06497_ net805 _01623_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08236_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__inv_2
XANTENNA__09966__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ net282 net490 vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nor2_1
XANTENNA__10905__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09267__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ top.DUT.register\[27\]\[12\] net777 net714 top.DUT.register\[30\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ _03223_ _03224_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12407__RESET_B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_189_Right_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06621__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ top.DUT.register\[6\]\[10\] net763 net673 top.DUT.register\[16\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_54_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ net154 net2121 net423 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07515__A _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Left_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ net1286 _04987_ _04979_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ clknet_leaf_91_clk _01293_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[35\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_178_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12701_ clknet_leaf_108_clk _00265_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13681_ clknet_leaf_94_clk _00007_ net993 vssd1 vssd1 vccd1 vccd1 top.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10893_ net1556 net176 net345 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ clknet_leaf_109_clk _00196_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08346__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10087__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ clknet_leaf_2_clk _00127_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11514_ _05349_ _05371_ _05361_ _05353_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ clknet_leaf_82_clk _00061_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramstore\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06860__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ _05289_ _05290_ _05272_ _05280_ _05281_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10815__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08081__A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ _05201_ _05226_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07404__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06612__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ net1423 net174 net398 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
X_13115_ clknet_leaf_56_clk _00679_ net1087 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13046_ clknet_leaf_2_clk _00610_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10258_ net1623 net172 net456 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__mux2_1
XANTENNA__12877__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10550__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10189_ net185 net1680 net411 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08808__X _03910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06679__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ net1130 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06420_ _01528_ _01530_ _01542_ _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__or4_4
XFILLER_0_57_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07891__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06351_ top.d_ready _01478_ _01481_ _01482_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or4_4
XFILLER_0_17_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09070_ _02588_ _02634_ _02684_ _03524_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or4_1
X_06282_ net1675 net875 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[26\] sky130_fd_sc_hd__and2_1
XANTENNA__07643__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08021_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__inv_2
XANTENNA__06851__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold702 top.DUT.register\[24\]\[6\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12571__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09087__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold713 top.DUT.register\[5\]\[15\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_1__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold724 top.DUT.register\[5\]\[2\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 top.DUT.register\[7\]\[22\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold746 top.DUT.register\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12500__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold757 top.DUT.register\[14\]\[4\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06603__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold768 top.DUT.register\[30\]\[7\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 top.DUT.register\[9\]\[27\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ net1550 net224 net429 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08923_ net286 _03289_ _03347_ net303 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o31a_1
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net474 _03942_ _03944_ net471 _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1004_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ top.DUT.register\[1\]\[19\] net657 net550 top.DUT.register\[24\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _03194_ _03206_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__nand2_1
XANTENNA__09305__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ top.DUT.register\[4\]\[1\] net769 net709 top.DUT.register\[9\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09856__B1 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07667_ top.DUT.register\[4\]\[0\] net564 net552 top.DUT.register\[7\]\[0\] _02793_
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout631_A _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06618_ top.DUT.register\[9\]\[28\] net709 net691 top.DUT.register\[3\]\[28\] _01744_
+ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ _01619_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07882__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ top.DUT.register\[23\]\[3\] net696 net685 top.DUT.register\[1\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XANTENNA__12207__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ net907 top.pc\[16\] _04382_ _04384_ top.testpc.en_latched vssd1 vssd1 vccd1
+ vccd1 _00097_ sky130_fd_sc_hd__o221a_1
X_06549_ top.DUT.register\[25\]\[30\] net623 net612 top.DUT.register\[14\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__a22o_1
XANTENNA__10983__X _05004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09268_ _04302_ _04306_ _04305_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08831__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__X _03572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ _02877_ net488 net481 _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09199_ top.pc\[8\] _04241_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nor2_1
XANTENNA__10635__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ net879 net880 _05098_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ net1338 net532 net525 _05068_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__a22o_1
X_10112_ net1601 net196 net461 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XANTENNA__09725__A _04718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ net914 net1304 net854 _05032_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a31o_1
XANTENNA__08347__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ net207 top.DUT.register\[5\]\[12\] net422 vssd1 vssd1 vccd1 vccd1 _00262_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08898__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 top.a1.row1\[2\] vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _01180_ vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 top.ramstore\[22\] vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 top.ramstore\[31\] vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 top.a1.data\[9\] vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _01169_ vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11990__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13802_ clknet_leaf_64_clk _01345_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11994_ _05862_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13733_ clknet_leaf_74_clk _01276_ net1089 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ _04629_ net849 vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nand2_4
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13664_ clknet_leaf_86_clk _01223_ net1007 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
X_10876_ top.DUT.register\[30\]\[6\] net245 net347 vssd1 vssd1 vccd1 vccd1 _01056_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07873__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12615_ clknet_leaf_26_clk _00179_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13595_ clknet_leaf_96_clk _01154_ net987 vssd1 vssd1 vccd1 vccd1 top.ramload\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07086__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__X _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07625__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ clknet_leaf_80_clk _00110_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[29\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_136_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06833__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10545__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ clknet_leaf_95_clk top.ru.next_FetchedInstr\[29\] net994 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[29\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_4 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11428_ top.a1.dataIn\[16\] _05295_ _05296_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08586__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ top.a1.dataIn\[27\] _05228_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09906__Y _04900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__D _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10280__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13029_ clknet_leaf_119_clk _00593_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_206_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1060 net1068 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
XANTENNA__07010__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1071 net1076 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_2
XANTENNA__13117__RESET_B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1093 net1097 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08570_ _02318_ net488 net486 _02319_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__a2bb2o_1
X_07521_ top.DUT.register\[23\]\[4\] net562 net637 top.DUT.register\[16\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10999__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07452_ top.DUT.register\[26\]\[6\] net621 _02570_ _02576_ _02578_ vssd1 vssd1 vccd1
+ vccd1 _02579_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06403_ top.DUT.register\[22\]\[30\] net751 net719 top.DUT.register\[2\]\[30\] _01524_
+ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07383_ top.DUT.register\[23\]\[7\] net696 _02502_ _02509_ vssd1 vssd1 vccd1 vccd1
+ _02510_ sky130_fd_sc_hd__a211o_1
X_09122_ net895 top.pc\[3\] vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or2_1
X_06334_ _01335_ _01460_ _01470_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__o21a_1
XANTENNA__07616__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08813__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _04106_ _04110_ _04111_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__and4_1
XFILLER_0_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06265_ net1302 net876 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[9\] sky130_fd_sc_hd__and2_1
XANTENNA__10455__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ top.DUT.register\[17\]\[31\] net645 net602 top.DUT.register\[10\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 top.DUT.register\[16\]\[19\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
X_06196_ net2261 _01419_ _01422_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[7\] sky130_fd_sc_hd__a21o_1
XFILLER_0_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold521 top.DUT.register\[25\]\[4\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold532 top.DUT.register\[23\]\[19\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold543 top.DUT.register\[30\]\[19\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 top.DUT.register\[24\]\[5\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 top.DUT.register\[4\]\[5\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 top.DUT.register\[23\]\[16\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 top.DUT.register\[27\]\[19\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 top.DUT.register\[4\]\[13\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06521__X _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ net162 net2077 net434 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout581_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net305 _04001_ _04002_ net273 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a211o_1
XANTENNA__10190__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10136__A0 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ top.pc\[28\] _04578_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__nand2_1
XANTENNA__07001__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07065__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08837_ _03916_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08768_ _03266_ _03269_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09280__A _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07719_ top.DUT.register\[11\]\[1\] net641 net609 top.DUT.register\[12\]\[1\] _02845_
+ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ net176 net2157 net381 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07855__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ net1426 net214 net452 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12400_ clknet_leaf_83_clk _00036_ net1013 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09279__X _04330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ clknet_leaf_40_clk _00944_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ net201 net2172 net387 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12331_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[1\]
+ top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12262_ top.lcd.cnt_20ms\[9\] top.lcd.cnt_20ms\[8\] _06081_ top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ net879 top.lcd.nextState\[4\] net892 net880 vssd1 vssd1 vccd1 vccd1 _05093_
+ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_186_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12193_ net1452 net846 net814 _06053_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__a22o_1
XANTENNA__08630__Y _03741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
X_11144_ net914 net1358 net853 _05058_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a31o_1
XANTENNA__07240__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06594__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ net91 net863 net826 net1241 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a22o_1
X_10026_ net154 net1836 net426 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_201_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _05825_ _05845_ _05752_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13716_ clknet_leaf_72_clk _01264_ net1096 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[13\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07846__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10928_ net169 net1295 net442 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09048__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ clknet_leaf_84_clk _01206_ net1015 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
X_10859_ net1633 net185 net351 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09599__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_167_Left_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ clknet_leaf_96_clk _01137_ net983 vssd1 vssd1 vccd1 vccd1 top.ramload\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06806__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ clknet_leaf_81_clk _00093_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11158__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__C1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13369__RESET_B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07584__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
Xfanout319 net321 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09740_ net833 _04343_ _04349_ net527 vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a2bb2o_1
X_06952_ _02077_ _02078_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__or2_2
.ends

